/* Machine-generated using LiteX gen */
module top(
	input clk100,
	input cpu_reset,
	output reg serial_tx,
	input serial_rx,
	input user_sw0,
	output oled_dc,
	output oled_res,
	output oled_sclk,
	output oled_sdin,
	output oled_vbat,
	output oled_vdd,
	output [14:0] ddram_a,
	output [2:0] ddram_ba,
	output ddram_ras_n,
	output ddram_cas_n,
	output ddram_we_n,
	output [1:0] ddram_dm,
	inout [15:0] ddram_dq,
	output [1:0] ddram_dqs_p,
	output [1:0] ddram_dqs_n,
	output ddram_clk_p,
	output ddram_clk_n,
	output ddram_cke,
	output ddram_odt,
	output ddram_reset_n,
	output reg spiflash_1x_cs_n,
	output reg spiflash_1x_mosi,
	input spiflash_1x_miso,
	output spiflash_1x_wp,
	output spiflash_1x_hold,
	output eth_clocks_tx,
	input eth_clocks_rx,
	output eth_rst_n,
	input eth_int_n,
	inout eth_mdio,
	output eth_mdc,
	input eth_rx_ctl,
	input [3:0] eth_rx_data,
	output eth_tx_ctl,
	output [3:0] eth_tx_data,
	input hdmi_in_clk_p,
	input hdmi_in_clk_n,
	input hdmi_in_data0_p,
	input hdmi_in_data0_n,
	input hdmi_in_data1_p,
	input hdmi_in_data1_n,
	input hdmi_in_data2_p,
	input hdmi_in_data2_n,
	input hdmi_in_scl,
	inout hdmi_in_sda,
	output hdmi_in_hpd_en,
	input hdmi_in_cec,
	output hdmi_in_txen,
	output hdmi_out_clk_p,
	output hdmi_out_clk_n,
	output hdmi_out_data0_p,
	output hdmi_out_data0_n,
	output hdmi_out_data1_p,
	output hdmi_out_data1_n,
	output hdmi_out_data2_p,
	output hdmi_out_data2_n,
	input hdmi_out_scl,
	input hdmi_out_sda,
	input hdmi_out_cec,
	input hdmi_out_hdp
);

wire [29:0] soc_videosoc_videosoc_ibus_adr;
wire [31:0] soc_videosoc_videosoc_ibus_dat_w;
wire [31:0] soc_videosoc_videosoc_ibus_dat_r;
wire [3:0] soc_videosoc_videosoc_ibus_sel;
wire soc_videosoc_videosoc_ibus_cyc;
wire soc_videosoc_videosoc_ibus_stb;
wire soc_videosoc_videosoc_ibus_ack;
wire soc_videosoc_videosoc_ibus_we;
wire [2:0] soc_videosoc_videosoc_ibus_cti;
wire [1:0] soc_videosoc_videosoc_ibus_bte;
wire soc_videosoc_videosoc_ibus_err;
wire [29:0] soc_videosoc_videosoc_dbus_adr;
wire [31:0] soc_videosoc_videosoc_dbus_dat_w;
wire [31:0] soc_videosoc_videosoc_dbus_dat_r;
wire [3:0] soc_videosoc_videosoc_dbus_sel;
wire soc_videosoc_videosoc_dbus_cyc;
wire soc_videosoc_videosoc_dbus_stb;
wire soc_videosoc_videosoc_dbus_ack;
wire soc_videosoc_videosoc_dbus_we;
wire [2:0] soc_videosoc_videosoc_dbus_cti;
wire [1:0] soc_videosoc_videosoc_dbus_bte;
wire soc_videosoc_videosoc_dbus_err;
reg [31:0] soc_videosoc_videosoc_interrupt = 32'd0;
wire [31:0] soc_videosoc_videosoc_i_adr_o;
wire [31:0] soc_videosoc_videosoc_d_adr_o;
wire [29:0] soc_videosoc_videosoc_rom_bus_adr;
wire [31:0] soc_videosoc_videosoc_rom_bus_dat_w;
wire [31:0] soc_videosoc_videosoc_rom_bus_dat_r;
wire [3:0] soc_videosoc_videosoc_rom_bus_sel;
wire soc_videosoc_videosoc_rom_bus_cyc;
wire soc_videosoc_videosoc_rom_bus_stb;
reg soc_videosoc_videosoc_rom_bus_ack = 1'd0;
wire soc_videosoc_videosoc_rom_bus_we;
wire [2:0] soc_videosoc_videosoc_rom_bus_cti;
wire [1:0] soc_videosoc_videosoc_rom_bus_bte;
reg soc_videosoc_videosoc_rom_bus_err = 1'd0;
wire [12:0] soc_videosoc_videosoc_rom_adr;
wire [31:0] soc_videosoc_videosoc_rom_dat_r;
wire [29:0] soc_videosoc_videosoc_sram_bus_adr;
wire [31:0] soc_videosoc_videosoc_sram_bus_dat_w;
wire [31:0] soc_videosoc_videosoc_sram_bus_dat_r;
wire [3:0] soc_videosoc_videosoc_sram_bus_sel;
wire soc_videosoc_videosoc_sram_bus_cyc;
wire soc_videosoc_videosoc_sram_bus_stb;
reg soc_videosoc_videosoc_sram_bus_ack = 1'd0;
wire soc_videosoc_videosoc_sram_bus_we;
wire [2:0] soc_videosoc_videosoc_sram_bus_cti;
wire [1:0] soc_videosoc_videosoc_sram_bus_bte;
reg soc_videosoc_videosoc_sram_bus_err = 1'd0;
wire [12:0] soc_videosoc_videosoc_sram_adr;
wire [31:0] soc_videosoc_videosoc_sram_dat_r;
reg [3:0] soc_videosoc_videosoc_sram_we = 4'd0;
wire [31:0] soc_videosoc_videosoc_sram_dat_w;
reg [13:0] soc_videosoc_videosoc_interface_adr = 14'd0;
reg soc_videosoc_videosoc_interface_we = 1'd0;
reg [7:0] soc_videosoc_videosoc_interface_dat_w = 8'd0;
wire [7:0] soc_videosoc_videosoc_interface_dat_r;
wire [29:0] soc_videosoc_videosoc_bus_wishbone_adr;
wire [31:0] soc_videosoc_videosoc_bus_wishbone_dat_w;
reg [31:0] soc_videosoc_videosoc_bus_wishbone_dat_r = 32'd0;
wire [3:0] soc_videosoc_videosoc_bus_wishbone_sel;
wire soc_videosoc_videosoc_bus_wishbone_cyc;
wire soc_videosoc_videosoc_bus_wishbone_stb;
reg soc_videosoc_videosoc_bus_wishbone_ack = 1'd0;
wire soc_videosoc_videosoc_bus_wishbone_we;
wire [2:0] soc_videosoc_videosoc_bus_wishbone_cti;
wire [1:0] soc_videosoc_videosoc_bus_wishbone_bte;
reg soc_videosoc_videosoc_bus_wishbone_err = 1'd0;
reg [1:0] soc_videosoc_videosoc_counter = 2'd0;
reg [31:0] soc_videosoc_videosoc_load_storage_full = 32'd0;
wire [31:0] soc_videosoc_videosoc_load_storage;
reg soc_videosoc_videosoc_load_re = 1'd0;
reg [31:0] soc_videosoc_videosoc_reload_storage_full = 32'd0;
wire [31:0] soc_videosoc_videosoc_reload_storage;
reg soc_videosoc_videosoc_reload_re = 1'd0;
reg soc_videosoc_videosoc_en_storage_full = 1'd0;
wire soc_videosoc_videosoc_en_storage;
reg soc_videosoc_videosoc_en_re = 1'd0;
wire soc_videosoc_videosoc_update_value_re;
wire soc_videosoc_videosoc_update_value_r;
reg soc_videosoc_videosoc_update_value_w = 1'd0;
reg [31:0] soc_videosoc_videosoc_value_status = 32'd0;
wire soc_videosoc_videosoc_irq;
wire soc_videosoc_videosoc_zero_status;
reg soc_videosoc_videosoc_zero_pending = 1'd0;
wire soc_videosoc_videosoc_zero_trigger;
reg soc_videosoc_videosoc_zero_clear = 1'd0;
reg soc_videosoc_videosoc_zero_old_trigger = 1'd0;
wire soc_videosoc_videosoc_eventmanager_status_re;
wire soc_videosoc_videosoc_eventmanager_status_r;
wire soc_videosoc_videosoc_eventmanager_status_w;
wire soc_videosoc_videosoc_eventmanager_pending_re;
wire soc_videosoc_videosoc_eventmanager_pending_r;
wire soc_videosoc_videosoc_eventmanager_pending_w;
reg soc_videosoc_videosoc_eventmanager_storage_full = 1'd0;
wire soc_videosoc_videosoc_eventmanager_storage;
reg soc_videosoc_videosoc_eventmanager_re = 1'd0;
reg [31:0] soc_videosoc_videosoc_value = 32'd0;
wire [29:0] soc_videosoc_interface0_wb_sdram_adr;
wire [31:0] soc_videosoc_interface0_wb_sdram_dat_w;
reg [31:0] soc_videosoc_interface0_wb_sdram_dat_r = 32'd0;
wire [3:0] soc_videosoc_interface0_wb_sdram_sel;
wire soc_videosoc_interface0_wb_sdram_cyc;
wire soc_videosoc_interface0_wb_sdram_stb;
reg soc_videosoc_interface0_wb_sdram_ack = 1'd0;
wire soc_videosoc_interface0_wb_sdram_we;
wire [2:0] soc_videosoc_interface0_wb_sdram_cti;
wire [1:0] soc_videosoc_interface0_wb_sdram_bte;
reg soc_videosoc_interface0_wb_sdram_err = 1'd0;
(* dont_touch = "true" *) wire sys_clk;
wire sys_rst;
wire sys4x_clk;
wire sys4x_dqs_clk;
wire clk200_clk;
wire clk200_rst;
wire clk100_clk;
wire clk100_rst;
wire soc_videosoc_pll_locked;
wire soc_videosoc_pll_fb;
wire soc_videosoc_pll_sys;
wire soc_videosoc_pll_sys4x;
wire soc_videosoc_pll_sys4x_dqs;
wire soc_videosoc_pll_clk200;
reg [3:0] soc_videosoc_reset_counter = 4'd15;
reg soc_videosoc_ic_reset = 1'd1;
wire soc_videosoc_rs232phyinterface0_sink_valid;
reg soc_videosoc_rs232phyinterface0_sink_ready = 1'd0;
wire soc_videosoc_rs232phyinterface0_sink_first;
wire soc_videosoc_rs232phyinterface0_sink_last;
wire [7:0] soc_videosoc_rs232phyinterface0_sink_payload_data;
reg soc_videosoc_rs232phyinterface0_source_valid = 1'd0;
wire soc_videosoc_rs232phyinterface0_source_ready;
reg soc_videosoc_rs232phyinterface0_source_first = 1'd0;
reg soc_videosoc_rs232phyinterface0_source_last = 1'd0;
reg [7:0] soc_videosoc_rs232phyinterface0_source_payload_data = 8'd0;
reg soc_videosoc_rs232phyinterface1_sink_valid = 1'd0;
reg soc_videosoc_rs232phyinterface1_sink_ready = 1'd0;
reg soc_videosoc_rs232phyinterface1_sink_first = 1'd0;
wire soc_videosoc_rs232phyinterface1_sink_last;
reg [7:0] soc_videosoc_rs232phyinterface1_sink_payload_data = 8'd0;
reg soc_videosoc_rs232phyinterface1_source_valid = 1'd0;
wire soc_videosoc_rs232phyinterface1_source_ready;
reg soc_videosoc_rs232phyinterface1_source_first = 1'd0;
reg soc_videosoc_rs232phyinterface1_source_last = 1'd0;
reg [7:0] soc_videosoc_rs232phyinterface1_source_payload_data = 8'd0;
wire soc_videosoc_uart_rxtx_re;
wire [7:0] soc_videosoc_uart_rxtx_r;
wire [7:0] soc_videosoc_uart_rxtx_w;
wire soc_videosoc_uart_txfull_status;
wire soc_videosoc_uart_rxempty_status;
wire soc_videosoc_uart_irq;
wire soc_videosoc_uart_tx_status;
reg soc_videosoc_uart_tx_pending = 1'd0;
wire soc_videosoc_uart_tx_trigger;
reg soc_videosoc_uart_tx_clear = 1'd0;
reg soc_videosoc_uart_tx_old_trigger = 1'd0;
wire soc_videosoc_uart_rx_status;
reg soc_videosoc_uart_rx_pending = 1'd0;
wire soc_videosoc_uart_rx_trigger;
reg soc_videosoc_uart_rx_clear = 1'd0;
reg soc_videosoc_uart_rx_old_trigger = 1'd0;
wire soc_videosoc_uart_status_re;
wire [1:0] soc_videosoc_uart_status_r;
reg [1:0] soc_videosoc_uart_status_w = 2'd0;
wire soc_videosoc_uart_pending_re;
wire [1:0] soc_videosoc_uart_pending_r;
reg [1:0] soc_videosoc_uart_pending_w = 2'd0;
reg [1:0] soc_videosoc_uart_storage_full = 2'd0;
wire [1:0] soc_videosoc_uart_storage;
reg soc_videosoc_uart_re = 1'd0;
wire soc_videosoc_uart_tx_fifo_sink_valid;
wire soc_videosoc_uart_tx_fifo_sink_ready;
reg soc_videosoc_uart_tx_fifo_sink_first = 1'd0;
reg soc_videosoc_uart_tx_fifo_sink_last = 1'd0;
wire [7:0] soc_videosoc_uart_tx_fifo_sink_payload_data;
wire soc_videosoc_uart_tx_fifo_source_valid;
wire soc_videosoc_uart_tx_fifo_source_ready;
wire soc_videosoc_uart_tx_fifo_source_first;
wire soc_videosoc_uart_tx_fifo_source_last;
wire [7:0] soc_videosoc_uart_tx_fifo_source_payload_data;
wire soc_videosoc_uart_tx_fifo_syncfifo_we;
wire soc_videosoc_uart_tx_fifo_syncfifo_writable;
wire soc_videosoc_uart_tx_fifo_syncfifo_re;
wire soc_videosoc_uart_tx_fifo_syncfifo_readable;
wire [9:0] soc_videosoc_uart_tx_fifo_syncfifo_din;
wire [9:0] soc_videosoc_uart_tx_fifo_syncfifo_dout;
reg [4:0] soc_videosoc_uart_tx_fifo_level = 5'd0;
reg soc_videosoc_uart_tx_fifo_replace = 1'd0;
reg [3:0] soc_videosoc_uart_tx_fifo_produce = 4'd0;
reg [3:0] soc_videosoc_uart_tx_fifo_consume = 4'd0;
reg [3:0] soc_videosoc_uart_tx_fifo_wrport_adr = 4'd0;
wire [9:0] soc_videosoc_uart_tx_fifo_wrport_dat_r;
wire soc_videosoc_uart_tx_fifo_wrport_we;
wire [9:0] soc_videosoc_uart_tx_fifo_wrport_dat_w;
wire soc_videosoc_uart_tx_fifo_do_read;
wire [3:0] soc_videosoc_uart_tx_fifo_rdport_adr;
wire [9:0] soc_videosoc_uart_tx_fifo_rdport_dat_r;
wire [7:0] soc_videosoc_uart_tx_fifo_fifo_in_payload_data;
wire soc_videosoc_uart_tx_fifo_fifo_in_first;
wire soc_videosoc_uart_tx_fifo_fifo_in_last;
wire [7:0] soc_videosoc_uart_tx_fifo_fifo_out_payload_data;
wire soc_videosoc_uart_tx_fifo_fifo_out_first;
wire soc_videosoc_uart_tx_fifo_fifo_out_last;
wire soc_videosoc_uart_rx_fifo_sink_valid;
wire soc_videosoc_uart_rx_fifo_sink_ready;
wire soc_videosoc_uart_rx_fifo_sink_first;
wire soc_videosoc_uart_rx_fifo_sink_last;
wire [7:0] soc_videosoc_uart_rx_fifo_sink_payload_data;
wire soc_videosoc_uart_rx_fifo_source_valid;
wire soc_videosoc_uart_rx_fifo_source_ready;
wire soc_videosoc_uart_rx_fifo_source_first;
wire soc_videosoc_uart_rx_fifo_source_last;
wire [7:0] soc_videosoc_uart_rx_fifo_source_payload_data;
wire soc_videosoc_uart_rx_fifo_syncfifo_we;
wire soc_videosoc_uart_rx_fifo_syncfifo_writable;
wire soc_videosoc_uart_rx_fifo_syncfifo_re;
wire soc_videosoc_uart_rx_fifo_syncfifo_readable;
wire [9:0] soc_videosoc_uart_rx_fifo_syncfifo_din;
wire [9:0] soc_videosoc_uart_rx_fifo_syncfifo_dout;
reg [4:0] soc_videosoc_uart_rx_fifo_level = 5'd0;
reg soc_videosoc_uart_rx_fifo_replace = 1'd0;
reg [3:0] soc_videosoc_uart_rx_fifo_produce = 4'd0;
reg [3:0] soc_videosoc_uart_rx_fifo_consume = 4'd0;
reg [3:0] soc_videosoc_uart_rx_fifo_wrport_adr = 4'd0;
wire [9:0] soc_videosoc_uart_rx_fifo_wrport_dat_r;
wire soc_videosoc_uart_rx_fifo_wrport_we;
wire [9:0] soc_videosoc_uart_rx_fifo_wrport_dat_w;
wire soc_videosoc_uart_rx_fifo_do_read;
wire [3:0] soc_videosoc_uart_rx_fifo_rdport_adr;
wire [9:0] soc_videosoc_uart_rx_fifo_rdport_dat_r;
wire [7:0] soc_videosoc_uart_rx_fifo_fifo_in_payload_data;
wire soc_videosoc_uart_rx_fifo_fifo_in_first;
wire soc_videosoc_uart_rx_fifo_fifo_in_last;
wire [7:0] soc_videosoc_uart_rx_fifo_fifo_out_payload_data;
wire soc_videosoc_uart_rx_fifo_fifo_out_first;
wire soc_videosoc_uart_rx_fifo_fifo_out_last;
wire [29:0] soc_videosoc_bridge_wishbone_adr;
wire [31:0] soc_videosoc_bridge_wishbone_dat_w;
wire [31:0] soc_videosoc_bridge_wishbone_dat_r;
wire [3:0] soc_videosoc_bridge_wishbone_sel;
reg soc_videosoc_bridge_wishbone_cyc = 1'd0;
reg soc_videosoc_bridge_wishbone_stb = 1'd0;
wire soc_videosoc_bridge_wishbone_ack;
reg soc_videosoc_bridge_wishbone_we = 1'd0;
reg [2:0] soc_videosoc_bridge_wishbone_cti = 3'd0;
reg [1:0] soc_videosoc_bridge_wishbone_bte = 2'd0;
wire soc_videosoc_bridge_wishbone_err;
reg [2:0] soc_videosoc_bridge_byte_counter = 3'd0;
reg soc_videosoc_bridge_byte_counter_reset = 1'd0;
reg soc_videosoc_bridge_byte_counter_ce = 1'd0;
reg [2:0] soc_videosoc_bridge_word_counter = 3'd0;
reg soc_videosoc_bridge_word_counter_reset = 1'd0;
reg soc_videosoc_bridge_word_counter_ce = 1'd0;
reg [7:0] soc_videosoc_bridge_cmd = 8'd0;
reg soc_videosoc_bridge_cmd_ce = 1'd0;
reg [7:0] soc_videosoc_bridge_length = 8'd0;
reg soc_videosoc_bridge_length_ce = 1'd0;
reg [31:0] soc_videosoc_bridge_address = 32'd0;
reg soc_videosoc_bridge_address_ce = 1'd0;
reg [31:0] soc_videosoc_bridge_data = 32'd0;
reg soc_videosoc_bridge_rx_data_ce = 1'd0;
reg soc_videosoc_bridge_tx_data_ce = 1'd0;
wire soc_videosoc_bridge_reset;
wire soc_videosoc_bridge_wait;
wire soc_videosoc_bridge_done;
reg [23:0] soc_videosoc_bridge_count = 24'd10000000;
reg soc_videosoc_bridge_is_ongoing = 1'd0;
reg [31:0] soc_videosoc_uart_phy_storage_full = 32'd4947802;
wire [31:0] soc_videosoc_uart_phy_storage;
reg soc_videosoc_uart_phy_re = 1'd0;
reg soc_videosoc_uart_phy_sink_valid = 1'd0;
reg soc_videosoc_uart_phy_sink_ready = 1'd0;
reg soc_videosoc_uart_phy_sink_first = 1'd0;
reg soc_videosoc_uart_phy_sink_last = 1'd0;
reg [7:0] soc_videosoc_uart_phy_sink_payload_data = 8'd0;
reg soc_videosoc_uart_phy_uart_clk_txen = 1'd0;
reg [31:0] soc_videosoc_uart_phy_phase_accumulator_tx = 32'd0;
reg [7:0] soc_videosoc_uart_phy_tx_reg = 8'd0;
reg [3:0] soc_videosoc_uart_phy_tx_bitcount = 4'd0;
reg soc_videosoc_uart_phy_tx_busy = 1'd0;
reg soc_videosoc_uart_phy_source_valid = 1'd0;
reg soc_videosoc_uart_phy_source_ready = 1'd0;
reg soc_videosoc_uart_phy_source_first = 1'd0;
reg soc_videosoc_uart_phy_source_last = 1'd0;
reg [7:0] soc_videosoc_uart_phy_source_payload_data = 8'd0;
reg soc_videosoc_uart_phy_uart_clk_rxen = 1'd0;
reg [31:0] soc_videosoc_uart_phy_phase_accumulator_rx = 32'd0;
wire soc_videosoc_uart_phy_rx;
reg soc_videosoc_uart_phy_rx_r = 1'd0;
reg [7:0] soc_videosoc_uart_phy_rx_reg = 8'd0;
reg [3:0] soc_videosoc_uart_phy_rx_bitcount = 4'd0;
reg soc_videosoc_uart_phy_rx_busy = 1'd0;
wire soc_videosoc_sel;
reg [56:0] soc_videosoc_info_dna_status = 57'd0;
wire soc_videosoc_info_dna_do;
reg [6:0] soc_videosoc_info_dna_cnt = 7'd0;
wire [159:0] soc_videosoc_info_git_status;
wire [63:0] soc_videosoc_info_platform_status;
wire [63:0] soc_videosoc_info_target_status;
reg [11:0] soc_videosoc_info_temperature_status = 12'd0;
reg [11:0] soc_videosoc_info_vccint_status = 12'd0;
reg [11:0] soc_videosoc_info_vccaux_status = 12'd0;
reg [11:0] soc_videosoc_info_vccbram_status = 12'd0;
wire [7:0] soc_videosoc_info_alarm;
wire soc_videosoc_info_ot;
wire soc_videosoc_info_busy;
wire [6:0] soc_videosoc_info_channel;
wire soc_videosoc_info_eoc;
wire soc_videosoc_info_eos;
wire [15:0] soc_videosoc_info_data;
wire soc_videosoc_info_drdy;
wire soc_videosoc_oled_spi_pads_cs_n;
reg soc_videosoc_oled_spi_pads_clk = 1'd0;
reg soc_videosoc_oled_spi_pads_mosi = 1'd0;
wire soc_videosoc_oled_spimaster_ctrl_re;
wire soc_videosoc_oled_spimaster_ctrl_r;
reg soc_videosoc_oled_spimaster_ctrl_w = 1'd0;
reg [7:0] soc_videosoc_oled_spimaster_length_storage_full = 8'd0;
wire [7:0] soc_videosoc_oled_spimaster_length_storage;
reg soc_videosoc_oled_spimaster_length_re = 1'd0;
wire soc_videosoc_oled_spimaster_status;
reg [7:0] soc_videosoc_oled_spimaster_mosi_storage_full = 8'd0;
wire [7:0] soc_videosoc_oled_spimaster_mosi_storage;
reg soc_videosoc_oled_spimaster_mosi_re = 1'd0;
reg soc_videosoc_oled_spimaster_irq = 1'd0;
wire soc_videosoc_oled_spimaster_start;
reg soc_videosoc_oled_spimaster_enable_cs = 1'd0;
reg soc_videosoc_oled_spimaster_enable_shift = 1'd0;
reg soc_videosoc_oled_spimaster_done = 1'd0;
reg [3:0] soc_videosoc_oled_spimaster_i = 4'd0;
wire soc_videosoc_oled_spimaster_set_clk;
wire soc_videosoc_oled_spimaster_clr_clk;
reg [7:0] soc_videosoc_oled_spimaster_cnt = 8'd0;
reg soc_videosoc_oled_spimaster_clr_cnt = 1'd0;
reg soc_videosoc_oled_spimaster_inc_cnt = 1'd0;
reg [7:0] soc_videosoc_oled_spimaster_sr_mosi = 8'd0;
reg soc_videosoc_oled_spimaster = 1'd0;
reg [3:0] soc_videosoc_oled_storage_full = 4'd0;
wire [3:0] soc_videosoc_oled_storage;
reg soc_videosoc_oled_re = 1'd0;
reg [1:0] soc_videosoc_ddrphy_storage_full = 2'd0;
wire [1:0] soc_videosoc_ddrphy_storage;
reg soc_videosoc_ddrphy_re = 1'd0;
wire soc_videosoc_ddrphy_rdly_dq_rst_re;
wire soc_videosoc_ddrphy_rdly_dq_rst_r;
reg soc_videosoc_ddrphy_rdly_dq_rst_w = 1'd0;
wire soc_videosoc_ddrphy_rdly_dq_inc_re;
wire soc_videosoc_ddrphy_rdly_dq_inc_r;
reg soc_videosoc_ddrphy_rdly_dq_inc_w = 1'd0;
wire soc_videosoc_ddrphy_rdly_dq_bitslip_re;
wire soc_videosoc_ddrphy_rdly_dq_bitslip_r;
reg soc_videosoc_ddrphy_rdly_dq_bitslip_w = 1'd0;
wire [14:0] soc_videosoc_ddrphy_dfi_p0_address;
wire [2:0] soc_videosoc_ddrphy_dfi_p0_bank;
wire soc_videosoc_ddrphy_dfi_p0_cas_n;
wire soc_videosoc_ddrphy_dfi_p0_cs_n;
wire soc_videosoc_ddrphy_dfi_p0_ras_n;
wire soc_videosoc_ddrphy_dfi_p0_we_n;
wire soc_videosoc_ddrphy_dfi_p0_cke;
wire soc_videosoc_ddrphy_dfi_p0_odt;
wire soc_videosoc_ddrphy_dfi_p0_reset_n;
wire [31:0] soc_videosoc_ddrphy_dfi_p0_wrdata;
wire soc_videosoc_ddrphy_dfi_p0_wrdata_en;
wire [3:0] soc_videosoc_ddrphy_dfi_p0_wrdata_mask;
wire soc_videosoc_ddrphy_dfi_p0_rddata_en;
wire [31:0] soc_videosoc_ddrphy_dfi_p0_rddata;
reg soc_videosoc_ddrphy_dfi_p0_rddata_valid = 1'd0;
wire [14:0] soc_videosoc_ddrphy_dfi_p1_address;
wire [2:0] soc_videosoc_ddrphy_dfi_p1_bank;
wire soc_videosoc_ddrphy_dfi_p1_cas_n;
wire soc_videosoc_ddrphy_dfi_p1_cs_n;
wire soc_videosoc_ddrphy_dfi_p1_ras_n;
wire soc_videosoc_ddrphy_dfi_p1_we_n;
wire soc_videosoc_ddrphy_dfi_p1_cke;
wire soc_videosoc_ddrphy_dfi_p1_odt;
wire soc_videosoc_ddrphy_dfi_p1_reset_n;
wire [31:0] soc_videosoc_ddrphy_dfi_p1_wrdata;
wire soc_videosoc_ddrphy_dfi_p1_wrdata_en;
wire [3:0] soc_videosoc_ddrphy_dfi_p1_wrdata_mask;
wire soc_videosoc_ddrphy_dfi_p1_rddata_en;
wire [31:0] soc_videosoc_ddrphy_dfi_p1_rddata;
reg soc_videosoc_ddrphy_dfi_p1_rddata_valid = 1'd0;
wire [14:0] soc_videosoc_ddrphy_dfi_p2_address;
wire [2:0] soc_videosoc_ddrphy_dfi_p2_bank;
wire soc_videosoc_ddrphy_dfi_p2_cas_n;
wire soc_videosoc_ddrphy_dfi_p2_cs_n;
wire soc_videosoc_ddrphy_dfi_p2_ras_n;
wire soc_videosoc_ddrphy_dfi_p2_we_n;
wire soc_videosoc_ddrphy_dfi_p2_cke;
wire soc_videosoc_ddrphy_dfi_p2_odt;
wire soc_videosoc_ddrphy_dfi_p2_reset_n;
wire [31:0] soc_videosoc_ddrphy_dfi_p2_wrdata;
wire soc_videosoc_ddrphy_dfi_p2_wrdata_en;
wire [3:0] soc_videosoc_ddrphy_dfi_p2_wrdata_mask;
wire soc_videosoc_ddrphy_dfi_p2_rddata_en;
wire [31:0] soc_videosoc_ddrphy_dfi_p2_rddata;
reg soc_videosoc_ddrphy_dfi_p2_rddata_valid = 1'd0;
wire [14:0] soc_videosoc_ddrphy_dfi_p3_address;
wire [2:0] soc_videosoc_ddrphy_dfi_p3_bank;
wire soc_videosoc_ddrphy_dfi_p3_cas_n;
wire soc_videosoc_ddrphy_dfi_p3_cs_n;
wire soc_videosoc_ddrphy_dfi_p3_ras_n;
wire soc_videosoc_ddrphy_dfi_p3_we_n;
wire soc_videosoc_ddrphy_dfi_p3_cke;
wire soc_videosoc_ddrphy_dfi_p3_odt;
wire soc_videosoc_ddrphy_dfi_p3_reset_n;
wire [31:0] soc_videosoc_ddrphy_dfi_p3_wrdata;
wire soc_videosoc_ddrphy_dfi_p3_wrdata_en;
wire [3:0] soc_videosoc_ddrphy_dfi_p3_wrdata_mask;
wire soc_videosoc_ddrphy_dfi_p3_rddata_en;
wire [31:0] soc_videosoc_ddrphy_dfi_p3_rddata;
reg soc_videosoc_ddrphy_dfi_p3_rddata_valid = 1'd0;
wire soc_videosoc_ddrphy_sd_clk_se;
reg soc_videosoc_ddrphy_oe_dqs = 1'd0;
reg [7:0] soc_videosoc_ddrphy_dqs_serdes_pattern = 8'd85;
wire soc_videosoc_ddrphy_dqs0;
wire soc_videosoc_ddrphy_dqs_t0;
wire soc_videosoc_ddrphy_dqs1;
wire soc_videosoc_ddrphy_dqs_t1;
reg soc_videosoc_ddrphy_oe_dq = 1'd0;
wire soc_videosoc_ddrphy_dq_o0;
wire soc_videosoc_ddrphy_dq_i_nodelay0;
wire soc_videosoc_ddrphy_dq_i_delayed0;
wire soc_videosoc_ddrphy_dq_t0;
wire soc_videosoc_ddrphy_dq_o1;
wire soc_videosoc_ddrphy_dq_i_nodelay1;
wire soc_videosoc_ddrphy_dq_i_delayed1;
wire soc_videosoc_ddrphy_dq_t1;
wire soc_videosoc_ddrphy_dq_o2;
wire soc_videosoc_ddrphy_dq_i_nodelay2;
wire soc_videosoc_ddrphy_dq_i_delayed2;
wire soc_videosoc_ddrphy_dq_t2;
wire soc_videosoc_ddrphy_dq_o3;
wire soc_videosoc_ddrphy_dq_i_nodelay3;
wire soc_videosoc_ddrphy_dq_i_delayed3;
wire soc_videosoc_ddrphy_dq_t3;
wire soc_videosoc_ddrphy_dq_o4;
wire soc_videosoc_ddrphy_dq_i_nodelay4;
wire soc_videosoc_ddrphy_dq_i_delayed4;
wire soc_videosoc_ddrphy_dq_t4;
wire soc_videosoc_ddrphy_dq_o5;
wire soc_videosoc_ddrphy_dq_i_nodelay5;
wire soc_videosoc_ddrphy_dq_i_delayed5;
wire soc_videosoc_ddrphy_dq_t5;
wire soc_videosoc_ddrphy_dq_o6;
wire soc_videosoc_ddrphy_dq_i_nodelay6;
wire soc_videosoc_ddrphy_dq_i_delayed6;
wire soc_videosoc_ddrphy_dq_t6;
wire soc_videosoc_ddrphy_dq_o7;
wire soc_videosoc_ddrphy_dq_i_nodelay7;
wire soc_videosoc_ddrphy_dq_i_delayed7;
wire soc_videosoc_ddrphy_dq_t7;
wire soc_videosoc_ddrphy_dq_o8;
wire soc_videosoc_ddrphy_dq_i_nodelay8;
wire soc_videosoc_ddrphy_dq_i_delayed8;
wire soc_videosoc_ddrphy_dq_t8;
wire soc_videosoc_ddrphy_dq_o9;
wire soc_videosoc_ddrphy_dq_i_nodelay9;
wire soc_videosoc_ddrphy_dq_i_delayed9;
wire soc_videosoc_ddrphy_dq_t9;
wire soc_videosoc_ddrphy_dq_o10;
wire soc_videosoc_ddrphy_dq_i_nodelay10;
wire soc_videosoc_ddrphy_dq_i_delayed10;
wire soc_videosoc_ddrphy_dq_t10;
wire soc_videosoc_ddrphy_dq_o11;
wire soc_videosoc_ddrphy_dq_i_nodelay11;
wire soc_videosoc_ddrphy_dq_i_delayed11;
wire soc_videosoc_ddrphy_dq_t11;
wire soc_videosoc_ddrphy_dq_o12;
wire soc_videosoc_ddrphy_dq_i_nodelay12;
wire soc_videosoc_ddrphy_dq_i_delayed12;
wire soc_videosoc_ddrphy_dq_t12;
wire soc_videosoc_ddrphy_dq_o13;
wire soc_videosoc_ddrphy_dq_i_nodelay13;
wire soc_videosoc_ddrphy_dq_i_delayed13;
wire soc_videosoc_ddrphy_dq_t13;
wire soc_videosoc_ddrphy_dq_o14;
wire soc_videosoc_ddrphy_dq_i_nodelay14;
wire soc_videosoc_ddrphy_dq_i_delayed14;
wire soc_videosoc_ddrphy_dq_t14;
wire soc_videosoc_ddrphy_dq_o15;
wire soc_videosoc_ddrphy_dq_i_nodelay15;
wire soc_videosoc_ddrphy_dq_i_delayed15;
wire soc_videosoc_ddrphy_dq_t15;
reg soc_videosoc_ddrphy_n_rddata_en0 = 1'd0;
reg soc_videosoc_ddrphy_n_rddata_en1 = 1'd0;
reg soc_videosoc_ddrphy_n_rddata_en2 = 1'd0;
reg soc_videosoc_ddrphy_n_rddata_en3 = 1'd0;
reg soc_videosoc_ddrphy_n_rddata_en4 = 1'd0;
wire soc_videosoc_ddrphy_oe;
reg [3:0] soc_videosoc_ddrphy_last_wrdata_en = 4'd0;
wire [14:0] soc_videosoc_sdram_inti_p0_address;
wire [2:0] soc_videosoc_sdram_inti_p0_bank;
reg soc_videosoc_sdram_inti_p0_cas_n = 1'd1;
reg soc_videosoc_sdram_inti_p0_cs_n = 1'd1;
reg soc_videosoc_sdram_inti_p0_ras_n = 1'd1;
reg soc_videosoc_sdram_inti_p0_we_n = 1'd1;
wire soc_videosoc_sdram_inti_p0_cke;
wire soc_videosoc_sdram_inti_p0_odt;
wire soc_videosoc_sdram_inti_p0_reset_n;
wire [31:0] soc_videosoc_sdram_inti_p0_wrdata;
wire soc_videosoc_sdram_inti_p0_wrdata_en;
wire [3:0] soc_videosoc_sdram_inti_p0_wrdata_mask;
wire soc_videosoc_sdram_inti_p0_rddata_en;
reg [31:0] soc_videosoc_sdram_inti_p0_rddata = 32'd0;
reg soc_videosoc_sdram_inti_p0_rddata_valid = 1'd0;
wire [14:0] soc_videosoc_sdram_inti_p1_address;
wire [2:0] soc_videosoc_sdram_inti_p1_bank;
reg soc_videosoc_sdram_inti_p1_cas_n = 1'd1;
reg soc_videosoc_sdram_inti_p1_cs_n = 1'd1;
reg soc_videosoc_sdram_inti_p1_ras_n = 1'd1;
reg soc_videosoc_sdram_inti_p1_we_n = 1'd1;
wire soc_videosoc_sdram_inti_p1_cke;
wire soc_videosoc_sdram_inti_p1_odt;
wire soc_videosoc_sdram_inti_p1_reset_n;
wire [31:0] soc_videosoc_sdram_inti_p1_wrdata;
wire soc_videosoc_sdram_inti_p1_wrdata_en;
wire [3:0] soc_videosoc_sdram_inti_p1_wrdata_mask;
wire soc_videosoc_sdram_inti_p1_rddata_en;
reg [31:0] soc_videosoc_sdram_inti_p1_rddata = 32'd0;
reg soc_videosoc_sdram_inti_p1_rddata_valid = 1'd0;
wire [14:0] soc_videosoc_sdram_inti_p2_address;
wire [2:0] soc_videosoc_sdram_inti_p2_bank;
reg soc_videosoc_sdram_inti_p2_cas_n = 1'd1;
reg soc_videosoc_sdram_inti_p2_cs_n = 1'd1;
reg soc_videosoc_sdram_inti_p2_ras_n = 1'd1;
reg soc_videosoc_sdram_inti_p2_we_n = 1'd1;
wire soc_videosoc_sdram_inti_p2_cke;
wire soc_videosoc_sdram_inti_p2_odt;
wire soc_videosoc_sdram_inti_p2_reset_n;
wire [31:0] soc_videosoc_sdram_inti_p2_wrdata;
wire soc_videosoc_sdram_inti_p2_wrdata_en;
wire [3:0] soc_videosoc_sdram_inti_p2_wrdata_mask;
wire soc_videosoc_sdram_inti_p2_rddata_en;
reg [31:0] soc_videosoc_sdram_inti_p2_rddata = 32'd0;
reg soc_videosoc_sdram_inti_p2_rddata_valid = 1'd0;
wire [14:0] soc_videosoc_sdram_inti_p3_address;
wire [2:0] soc_videosoc_sdram_inti_p3_bank;
reg soc_videosoc_sdram_inti_p3_cas_n = 1'd1;
reg soc_videosoc_sdram_inti_p3_cs_n = 1'd1;
reg soc_videosoc_sdram_inti_p3_ras_n = 1'd1;
reg soc_videosoc_sdram_inti_p3_we_n = 1'd1;
wire soc_videosoc_sdram_inti_p3_cke;
wire soc_videosoc_sdram_inti_p3_odt;
wire soc_videosoc_sdram_inti_p3_reset_n;
wire [31:0] soc_videosoc_sdram_inti_p3_wrdata;
wire soc_videosoc_sdram_inti_p3_wrdata_en;
wire [3:0] soc_videosoc_sdram_inti_p3_wrdata_mask;
wire soc_videosoc_sdram_inti_p3_rddata_en;
reg [31:0] soc_videosoc_sdram_inti_p3_rddata = 32'd0;
reg soc_videosoc_sdram_inti_p3_rddata_valid = 1'd0;
wire [14:0] soc_videosoc_sdram_slave_p0_address;
wire [2:0] soc_videosoc_sdram_slave_p0_bank;
wire soc_videosoc_sdram_slave_p0_cas_n;
wire soc_videosoc_sdram_slave_p0_cs_n;
wire soc_videosoc_sdram_slave_p0_ras_n;
wire soc_videosoc_sdram_slave_p0_we_n;
wire soc_videosoc_sdram_slave_p0_cke;
wire soc_videosoc_sdram_slave_p0_odt;
wire soc_videosoc_sdram_slave_p0_reset_n;
wire [31:0] soc_videosoc_sdram_slave_p0_wrdata;
wire soc_videosoc_sdram_slave_p0_wrdata_en;
wire [3:0] soc_videosoc_sdram_slave_p0_wrdata_mask;
wire soc_videosoc_sdram_slave_p0_rddata_en;
reg [31:0] soc_videosoc_sdram_slave_p0_rddata = 32'd0;
reg soc_videosoc_sdram_slave_p0_rddata_valid = 1'd0;
wire [14:0] soc_videosoc_sdram_slave_p1_address;
wire [2:0] soc_videosoc_sdram_slave_p1_bank;
wire soc_videosoc_sdram_slave_p1_cas_n;
wire soc_videosoc_sdram_slave_p1_cs_n;
wire soc_videosoc_sdram_slave_p1_ras_n;
wire soc_videosoc_sdram_slave_p1_we_n;
wire soc_videosoc_sdram_slave_p1_cke;
wire soc_videosoc_sdram_slave_p1_odt;
wire soc_videosoc_sdram_slave_p1_reset_n;
wire [31:0] soc_videosoc_sdram_slave_p1_wrdata;
wire soc_videosoc_sdram_slave_p1_wrdata_en;
wire [3:0] soc_videosoc_sdram_slave_p1_wrdata_mask;
wire soc_videosoc_sdram_slave_p1_rddata_en;
reg [31:0] soc_videosoc_sdram_slave_p1_rddata = 32'd0;
reg soc_videosoc_sdram_slave_p1_rddata_valid = 1'd0;
wire [14:0] soc_videosoc_sdram_slave_p2_address;
wire [2:0] soc_videosoc_sdram_slave_p2_bank;
wire soc_videosoc_sdram_slave_p2_cas_n;
wire soc_videosoc_sdram_slave_p2_cs_n;
wire soc_videosoc_sdram_slave_p2_ras_n;
wire soc_videosoc_sdram_slave_p2_we_n;
wire soc_videosoc_sdram_slave_p2_cke;
wire soc_videosoc_sdram_slave_p2_odt;
wire soc_videosoc_sdram_slave_p2_reset_n;
wire [31:0] soc_videosoc_sdram_slave_p2_wrdata;
wire soc_videosoc_sdram_slave_p2_wrdata_en;
wire [3:0] soc_videosoc_sdram_slave_p2_wrdata_mask;
wire soc_videosoc_sdram_slave_p2_rddata_en;
reg [31:0] soc_videosoc_sdram_slave_p2_rddata = 32'd0;
reg soc_videosoc_sdram_slave_p2_rddata_valid = 1'd0;
wire [14:0] soc_videosoc_sdram_slave_p3_address;
wire [2:0] soc_videosoc_sdram_slave_p3_bank;
wire soc_videosoc_sdram_slave_p3_cas_n;
wire soc_videosoc_sdram_slave_p3_cs_n;
wire soc_videosoc_sdram_slave_p3_ras_n;
wire soc_videosoc_sdram_slave_p3_we_n;
wire soc_videosoc_sdram_slave_p3_cke;
wire soc_videosoc_sdram_slave_p3_odt;
wire soc_videosoc_sdram_slave_p3_reset_n;
wire [31:0] soc_videosoc_sdram_slave_p3_wrdata;
wire soc_videosoc_sdram_slave_p3_wrdata_en;
wire [3:0] soc_videosoc_sdram_slave_p3_wrdata_mask;
wire soc_videosoc_sdram_slave_p3_rddata_en;
reg [31:0] soc_videosoc_sdram_slave_p3_rddata = 32'd0;
reg soc_videosoc_sdram_slave_p3_rddata_valid = 1'd0;
reg [14:0] soc_videosoc_sdram_master_p0_address = 15'd0;
reg [2:0] soc_videosoc_sdram_master_p0_bank = 3'd0;
reg soc_videosoc_sdram_master_p0_cas_n = 1'd1;
reg soc_videosoc_sdram_master_p0_cs_n = 1'd1;
reg soc_videosoc_sdram_master_p0_ras_n = 1'd1;
reg soc_videosoc_sdram_master_p0_we_n = 1'd1;
reg soc_videosoc_sdram_master_p0_cke = 1'd0;
reg soc_videosoc_sdram_master_p0_odt = 1'd0;
reg soc_videosoc_sdram_master_p0_reset_n = 1'd0;
reg [31:0] soc_videosoc_sdram_master_p0_wrdata = 32'd0;
reg soc_videosoc_sdram_master_p0_wrdata_en = 1'd0;
reg [3:0] soc_videosoc_sdram_master_p0_wrdata_mask = 4'd0;
reg soc_videosoc_sdram_master_p0_rddata_en = 1'd0;
wire [31:0] soc_videosoc_sdram_master_p0_rddata;
wire soc_videosoc_sdram_master_p0_rddata_valid;
reg [14:0] soc_videosoc_sdram_master_p1_address = 15'd0;
reg [2:0] soc_videosoc_sdram_master_p1_bank = 3'd0;
reg soc_videosoc_sdram_master_p1_cas_n = 1'd1;
reg soc_videosoc_sdram_master_p1_cs_n = 1'd1;
reg soc_videosoc_sdram_master_p1_ras_n = 1'd1;
reg soc_videosoc_sdram_master_p1_we_n = 1'd1;
reg soc_videosoc_sdram_master_p1_cke = 1'd0;
reg soc_videosoc_sdram_master_p1_odt = 1'd0;
reg soc_videosoc_sdram_master_p1_reset_n = 1'd0;
reg [31:0] soc_videosoc_sdram_master_p1_wrdata = 32'd0;
reg soc_videosoc_sdram_master_p1_wrdata_en = 1'd0;
reg [3:0] soc_videosoc_sdram_master_p1_wrdata_mask = 4'd0;
reg soc_videosoc_sdram_master_p1_rddata_en = 1'd0;
wire [31:0] soc_videosoc_sdram_master_p1_rddata;
wire soc_videosoc_sdram_master_p1_rddata_valid;
reg [14:0] soc_videosoc_sdram_master_p2_address = 15'd0;
reg [2:0] soc_videosoc_sdram_master_p2_bank = 3'd0;
reg soc_videosoc_sdram_master_p2_cas_n = 1'd1;
reg soc_videosoc_sdram_master_p2_cs_n = 1'd1;
reg soc_videosoc_sdram_master_p2_ras_n = 1'd1;
reg soc_videosoc_sdram_master_p2_we_n = 1'd1;
reg soc_videosoc_sdram_master_p2_cke = 1'd0;
reg soc_videosoc_sdram_master_p2_odt = 1'd0;
reg soc_videosoc_sdram_master_p2_reset_n = 1'd0;
reg [31:0] soc_videosoc_sdram_master_p2_wrdata = 32'd0;
reg soc_videosoc_sdram_master_p2_wrdata_en = 1'd0;
reg [3:0] soc_videosoc_sdram_master_p2_wrdata_mask = 4'd0;
reg soc_videosoc_sdram_master_p2_rddata_en = 1'd0;
wire [31:0] soc_videosoc_sdram_master_p2_rddata;
wire soc_videosoc_sdram_master_p2_rddata_valid;
reg [14:0] soc_videosoc_sdram_master_p3_address = 15'd0;
reg [2:0] soc_videosoc_sdram_master_p3_bank = 3'd0;
reg soc_videosoc_sdram_master_p3_cas_n = 1'd1;
reg soc_videosoc_sdram_master_p3_cs_n = 1'd1;
reg soc_videosoc_sdram_master_p3_ras_n = 1'd1;
reg soc_videosoc_sdram_master_p3_we_n = 1'd1;
reg soc_videosoc_sdram_master_p3_cke = 1'd0;
reg soc_videosoc_sdram_master_p3_odt = 1'd0;
reg soc_videosoc_sdram_master_p3_reset_n = 1'd0;
reg [31:0] soc_videosoc_sdram_master_p3_wrdata = 32'd0;
reg soc_videosoc_sdram_master_p3_wrdata_en = 1'd0;
reg [3:0] soc_videosoc_sdram_master_p3_wrdata_mask = 4'd0;
reg soc_videosoc_sdram_master_p3_rddata_en = 1'd0;
wire [31:0] soc_videosoc_sdram_master_p3_rddata;
wire soc_videosoc_sdram_master_p3_rddata_valid;
reg [3:0] soc_videosoc_sdram_storage_full = 4'd0;
wire [3:0] soc_videosoc_sdram_storage;
reg soc_videosoc_sdram_re = 1'd0;
reg [5:0] soc_videosoc_sdram_phaseinjector0_command_storage_full = 6'd0;
wire [5:0] soc_videosoc_sdram_phaseinjector0_command_storage;
reg soc_videosoc_sdram_phaseinjector0_command_re = 1'd0;
wire soc_videosoc_sdram_phaseinjector0_command_issue_re;
wire soc_videosoc_sdram_phaseinjector0_command_issue_r;
reg soc_videosoc_sdram_phaseinjector0_command_issue_w = 1'd0;
reg [14:0] soc_videosoc_sdram_phaseinjector0_address_storage_full = 15'd0;
wire [14:0] soc_videosoc_sdram_phaseinjector0_address_storage;
reg soc_videosoc_sdram_phaseinjector0_address_re = 1'd0;
reg [2:0] soc_videosoc_sdram_phaseinjector0_baddress_storage_full = 3'd0;
wire [2:0] soc_videosoc_sdram_phaseinjector0_baddress_storage;
reg soc_videosoc_sdram_phaseinjector0_baddress_re = 1'd0;
reg [31:0] soc_videosoc_sdram_phaseinjector0_wrdata_storage_full = 32'd0;
wire [31:0] soc_videosoc_sdram_phaseinjector0_wrdata_storage;
reg soc_videosoc_sdram_phaseinjector0_wrdata_re = 1'd0;
reg [31:0] soc_videosoc_sdram_phaseinjector0_status = 32'd0;
reg [5:0] soc_videosoc_sdram_phaseinjector1_command_storage_full = 6'd0;
wire [5:0] soc_videosoc_sdram_phaseinjector1_command_storage;
reg soc_videosoc_sdram_phaseinjector1_command_re = 1'd0;
wire soc_videosoc_sdram_phaseinjector1_command_issue_re;
wire soc_videosoc_sdram_phaseinjector1_command_issue_r;
reg soc_videosoc_sdram_phaseinjector1_command_issue_w = 1'd0;
reg [14:0] soc_videosoc_sdram_phaseinjector1_address_storage_full = 15'd0;
wire [14:0] soc_videosoc_sdram_phaseinjector1_address_storage;
reg soc_videosoc_sdram_phaseinjector1_address_re = 1'd0;
reg [2:0] soc_videosoc_sdram_phaseinjector1_baddress_storage_full = 3'd0;
wire [2:0] soc_videosoc_sdram_phaseinjector1_baddress_storage;
reg soc_videosoc_sdram_phaseinjector1_baddress_re = 1'd0;
reg [31:0] soc_videosoc_sdram_phaseinjector1_wrdata_storage_full = 32'd0;
wire [31:0] soc_videosoc_sdram_phaseinjector1_wrdata_storage;
reg soc_videosoc_sdram_phaseinjector1_wrdata_re = 1'd0;
reg [31:0] soc_videosoc_sdram_phaseinjector1_status = 32'd0;
reg [5:0] soc_videosoc_sdram_phaseinjector2_command_storage_full = 6'd0;
wire [5:0] soc_videosoc_sdram_phaseinjector2_command_storage;
reg soc_videosoc_sdram_phaseinjector2_command_re = 1'd0;
wire soc_videosoc_sdram_phaseinjector2_command_issue_re;
wire soc_videosoc_sdram_phaseinjector2_command_issue_r;
reg soc_videosoc_sdram_phaseinjector2_command_issue_w = 1'd0;
reg [14:0] soc_videosoc_sdram_phaseinjector2_address_storage_full = 15'd0;
wire [14:0] soc_videosoc_sdram_phaseinjector2_address_storage;
reg soc_videosoc_sdram_phaseinjector2_address_re = 1'd0;
reg [2:0] soc_videosoc_sdram_phaseinjector2_baddress_storage_full = 3'd0;
wire [2:0] soc_videosoc_sdram_phaseinjector2_baddress_storage;
reg soc_videosoc_sdram_phaseinjector2_baddress_re = 1'd0;
reg [31:0] soc_videosoc_sdram_phaseinjector2_wrdata_storage_full = 32'd0;
wire [31:0] soc_videosoc_sdram_phaseinjector2_wrdata_storage;
reg soc_videosoc_sdram_phaseinjector2_wrdata_re = 1'd0;
reg [31:0] soc_videosoc_sdram_phaseinjector2_status = 32'd0;
reg [5:0] soc_videosoc_sdram_phaseinjector3_command_storage_full = 6'd0;
wire [5:0] soc_videosoc_sdram_phaseinjector3_command_storage;
reg soc_videosoc_sdram_phaseinjector3_command_re = 1'd0;
wire soc_videosoc_sdram_phaseinjector3_command_issue_re;
wire soc_videosoc_sdram_phaseinjector3_command_issue_r;
reg soc_videosoc_sdram_phaseinjector3_command_issue_w = 1'd0;
reg [14:0] soc_videosoc_sdram_phaseinjector3_address_storage_full = 15'd0;
wire [14:0] soc_videosoc_sdram_phaseinjector3_address_storage;
reg soc_videosoc_sdram_phaseinjector3_address_re = 1'd0;
reg [2:0] soc_videosoc_sdram_phaseinjector3_baddress_storage_full = 3'd0;
wire [2:0] soc_videosoc_sdram_phaseinjector3_baddress_storage;
reg soc_videosoc_sdram_phaseinjector3_baddress_re = 1'd0;
reg [31:0] soc_videosoc_sdram_phaseinjector3_wrdata_storage_full = 32'd0;
wire [31:0] soc_videosoc_sdram_phaseinjector3_wrdata_storage;
reg soc_videosoc_sdram_phaseinjector3_wrdata_re = 1'd0;
reg [31:0] soc_videosoc_sdram_phaseinjector3_status = 32'd0;
reg [14:0] soc_videosoc_sdram_dfi_p0_address = 15'd0;
reg [2:0] soc_videosoc_sdram_dfi_p0_bank = 3'd0;
reg soc_videosoc_sdram_dfi_p0_cas_n = 1'd1;
wire soc_videosoc_sdram_dfi_p0_cs_n;
reg soc_videosoc_sdram_dfi_p0_ras_n = 1'd1;
reg soc_videosoc_sdram_dfi_p0_we_n = 1'd1;
wire soc_videosoc_sdram_dfi_p0_cke;
wire soc_videosoc_sdram_dfi_p0_odt;
wire soc_videosoc_sdram_dfi_p0_reset_n;
wire [31:0] soc_videosoc_sdram_dfi_p0_wrdata;
reg soc_videosoc_sdram_dfi_p0_wrdata_en = 1'd0;
wire [3:0] soc_videosoc_sdram_dfi_p0_wrdata_mask;
reg soc_videosoc_sdram_dfi_p0_rddata_en = 1'd0;
wire [31:0] soc_videosoc_sdram_dfi_p0_rddata;
wire soc_videosoc_sdram_dfi_p0_rddata_valid;
reg [14:0] soc_videosoc_sdram_dfi_p1_address = 15'd0;
reg [2:0] soc_videosoc_sdram_dfi_p1_bank = 3'd0;
reg soc_videosoc_sdram_dfi_p1_cas_n = 1'd1;
wire soc_videosoc_sdram_dfi_p1_cs_n;
reg soc_videosoc_sdram_dfi_p1_ras_n = 1'd1;
reg soc_videosoc_sdram_dfi_p1_we_n = 1'd1;
wire soc_videosoc_sdram_dfi_p1_cke;
wire soc_videosoc_sdram_dfi_p1_odt;
wire soc_videosoc_sdram_dfi_p1_reset_n;
wire [31:0] soc_videosoc_sdram_dfi_p1_wrdata;
reg soc_videosoc_sdram_dfi_p1_wrdata_en = 1'd0;
wire [3:0] soc_videosoc_sdram_dfi_p1_wrdata_mask;
reg soc_videosoc_sdram_dfi_p1_rddata_en = 1'd0;
wire [31:0] soc_videosoc_sdram_dfi_p1_rddata;
wire soc_videosoc_sdram_dfi_p1_rddata_valid;
reg [14:0] soc_videosoc_sdram_dfi_p2_address = 15'd0;
reg [2:0] soc_videosoc_sdram_dfi_p2_bank = 3'd0;
reg soc_videosoc_sdram_dfi_p2_cas_n = 1'd1;
wire soc_videosoc_sdram_dfi_p2_cs_n;
reg soc_videosoc_sdram_dfi_p2_ras_n = 1'd1;
reg soc_videosoc_sdram_dfi_p2_we_n = 1'd1;
wire soc_videosoc_sdram_dfi_p2_cke;
wire soc_videosoc_sdram_dfi_p2_odt;
wire soc_videosoc_sdram_dfi_p2_reset_n;
wire [31:0] soc_videosoc_sdram_dfi_p2_wrdata;
reg soc_videosoc_sdram_dfi_p2_wrdata_en = 1'd0;
wire [3:0] soc_videosoc_sdram_dfi_p2_wrdata_mask;
reg soc_videosoc_sdram_dfi_p2_rddata_en = 1'd0;
wire [31:0] soc_videosoc_sdram_dfi_p2_rddata;
wire soc_videosoc_sdram_dfi_p2_rddata_valid;
reg [14:0] soc_videosoc_sdram_dfi_p3_address = 15'd0;
reg [2:0] soc_videosoc_sdram_dfi_p3_bank = 3'd0;
reg soc_videosoc_sdram_dfi_p3_cas_n = 1'd1;
wire soc_videosoc_sdram_dfi_p3_cs_n;
reg soc_videosoc_sdram_dfi_p3_ras_n = 1'd1;
reg soc_videosoc_sdram_dfi_p3_we_n = 1'd1;
wire soc_videosoc_sdram_dfi_p3_cke;
wire soc_videosoc_sdram_dfi_p3_odt;
wire soc_videosoc_sdram_dfi_p3_reset_n;
wire [31:0] soc_videosoc_sdram_dfi_p3_wrdata;
reg soc_videosoc_sdram_dfi_p3_wrdata_en = 1'd0;
wire [3:0] soc_videosoc_sdram_dfi_p3_wrdata_mask;
reg soc_videosoc_sdram_dfi_p3_rddata_en = 1'd0;
wire [31:0] soc_videosoc_sdram_dfi_p3_rddata;
wire soc_videosoc_sdram_dfi_p3_rddata_valid;
wire soc_videosoc_sdram_interface_bank0_valid;
wire soc_videosoc_sdram_interface_bank0_ready;
wire soc_videosoc_sdram_interface_bank0_we;
wire [21:0] soc_videosoc_sdram_interface_bank0_adr;
wire soc_videosoc_sdram_interface_bank0_lock;
wire soc_videosoc_sdram_interface_bank0_wdata_ready;
wire soc_videosoc_sdram_interface_bank0_rdata_valid;
wire soc_videosoc_sdram_interface_bank1_valid;
wire soc_videosoc_sdram_interface_bank1_ready;
wire soc_videosoc_sdram_interface_bank1_we;
wire [21:0] soc_videosoc_sdram_interface_bank1_adr;
wire soc_videosoc_sdram_interface_bank1_lock;
wire soc_videosoc_sdram_interface_bank1_wdata_ready;
wire soc_videosoc_sdram_interface_bank1_rdata_valid;
wire soc_videosoc_sdram_interface_bank2_valid;
wire soc_videosoc_sdram_interface_bank2_ready;
wire soc_videosoc_sdram_interface_bank2_we;
wire [21:0] soc_videosoc_sdram_interface_bank2_adr;
wire soc_videosoc_sdram_interface_bank2_lock;
wire soc_videosoc_sdram_interface_bank2_wdata_ready;
wire soc_videosoc_sdram_interface_bank2_rdata_valid;
wire soc_videosoc_sdram_interface_bank3_valid;
wire soc_videosoc_sdram_interface_bank3_ready;
wire soc_videosoc_sdram_interface_bank3_we;
wire [21:0] soc_videosoc_sdram_interface_bank3_adr;
wire soc_videosoc_sdram_interface_bank3_lock;
wire soc_videosoc_sdram_interface_bank3_wdata_ready;
wire soc_videosoc_sdram_interface_bank3_rdata_valid;
wire soc_videosoc_sdram_interface_bank4_valid;
wire soc_videosoc_sdram_interface_bank4_ready;
wire soc_videosoc_sdram_interface_bank4_we;
wire [21:0] soc_videosoc_sdram_interface_bank4_adr;
wire soc_videosoc_sdram_interface_bank4_lock;
wire soc_videosoc_sdram_interface_bank4_wdata_ready;
wire soc_videosoc_sdram_interface_bank4_rdata_valid;
wire soc_videosoc_sdram_interface_bank5_valid;
wire soc_videosoc_sdram_interface_bank5_ready;
wire soc_videosoc_sdram_interface_bank5_we;
wire [21:0] soc_videosoc_sdram_interface_bank5_adr;
wire soc_videosoc_sdram_interface_bank5_lock;
wire soc_videosoc_sdram_interface_bank5_wdata_ready;
wire soc_videosoc_sdram_interface_bank5_rdata_valid;
wire soc_videosoc_sdram_interface_bank6_valid;
wire soc_videosoc_sdram_interface_bank6_ready;
wire soc_videosoc_sdram_interface_bank6_we;
wire [21:0] soc_videosoc_sdram_interface_bank6_adr;
wire soc_videosoc_sdram_interface_bank6_lock;
wire soc_videosoc_sdram_interface_bank6_wdata_ready;
wire soc_videosoc_sdram_interface_bank6_rdata_valid;
wire soc_videosoc_sdram_interface_bank7_valid;
wire soc_videosoc_sdram_interface_bank7_ready;
wire soc_videosoc_sdram_interface_bank7_we;
wire [21:0] soc_videosoc_sdram_interface_bank7_adr;
wire soc_videosoc_sdram_interface_bank7_lock;
wire soc_videosoc_sdram_interface_bank7_wdata_ready;
wire soc_videosoc_sdram_interface_bank7_rdata_valid;
reg [127:0] soc_videosoc_sdram_interface_wdata = 128'd0;
reg [15:0] soc_videosoc_sdram_interface_wdata_we = 16'd0;
wire [127:0] soc_videosoc_sdram_interface_rdata;
reg soc_videosoc_sdram_cmd_valid = 1'd0;
reg soc_videosoc_sdram_cmd_ready = 1'd0;
reg soc_videosoc_sdram_cmd_last = 1'd0;
reg [14:0] soc_videosoc_sdram_cmd_payload_a = 15'd0;
reg [2:0] soc_videosoc_sdram_cmd_payload_ba = 3'd0;
reg soc_videosoc_sdram_cmd_payload_cas = 1'd0;
reg soc_videosoc_sdram_cmd_payload_ras = 1'd0;
reg soc_videosoc_sdram_cmd_payload_we = 1'd0;
reg soc_videosoc_sdram_cmd_payload_is_read = 1'd0;
reg soc_videosoc_sdram_cmd_payload_is_write = 1'd0;
reg soc_videosoc_sdram_seq_start = 1'd0;
reg soc_videosoc_sdram_seq_done = 1'd0;
reg [4:0] soc_videosoc_sdram_counter = 5'd0;
wire soc_videosoc_sdram_wait;
wire soc_videosoc_sdram_done;
reg [9:0] soc_videosoc_sdram_count = 10'd782;
wire soc_videosoc_sdram_bankmachine0_req_valid;
wire soc_videosoc_sdram_bankmachine0_req_ready;
wire soc_videosoc_sdram_bankmachine0_req_we;
wire [21:0] soc_videosoc_sdram_bankmachine0_req_adr;
wire soc_videosoc_sdram_bankmachine0_req_lock;
reg soc_videosoc_sdram_bankmachine0_req_wdata_ready = 1'd0;
reg soc_videosoc_sdram_bankmachine0_req_rdata_valid = 1'd0;
wire soc_videosoc_sdram_bankmachine0_refresh_req;
reg soc_videosoc_sdram_bankmachine0_refresh_gnt = 1'd0;
reg soc_videosoc_sdram_bankmachine0_cmd_valid = 1'd0;
reg soc_videosoc_sdram_bankmachine0_cmd_ready = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine0_cmd_payload_a = 15'd0;
wire [2:0] soc_videosoc_sdram_bankmachine0_cmd_payload_ba;
reg soc_videosoc_sdram_bankmachine0_cmd_payload_cas = 1'd0;
reg soc_videosoc_sdram_bankmachine0_cmd_payload_ras = 1'd0;
reg soc_videosoc_sdram_bankmachine0_cmd_payload_we = 1'd0;
reg soc_videosoc_sdram_bankmachine0_cmd_payload_is_cmd = 1'd0;
reg soc_videosoc_sdram_bankmachine0_cmd_payload_is_read = 1'd0;
reg soc_videosoc_sdram_bankmachine0_cmd_payload_is_write = 1'd0;
wire soc_videosoc_sdram_bankmachine0_sink_valid;
wire soc_videosoc_sdram_bankmachine0_sink_ready;
reg soc_videosoc_sdram_bankmachine0_sink_first = 1'd0;
reg soc_videosoc_sdram_bankmachine0_sink_last = 1'd0;
wire soc_videosoc_sdram_bankmachine0_sink_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine0_sink_payload_adr;
wire soc_videosoc_sdram_bankmachine0_source_valid;
wire soc_videosoc_sdram_bankmachine0_source_ready;
wire soc_videosoc_sdram_bankmachine0_source_first;
wire soc_videosoc_sdram_bankmachine0_source_last;
wire soc_videosoc_sdram_bankmachine0_source_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine0_source_payload_adr;
wire soc_videosoc_sdram_bankmachine0_syncfifo0_we;
wire soc_videosoc_sdram_bankmachine0_syncfifo0_writable;
wire soc_videosoc_sdram_bankmachine0_syncfifo0_re;
wire soc_videosoc_sdram_bankmachine0_syncfifo0_readable;
wire [24:0] soc_videosoc_sdram_bankmachine0_syncfifo0_din;
wire [24:0] soc_videosoc_sdram_bankmachine0_syncfifo0_dout;
reg [3:0] soc_videosoc_sdram_bankmachine0_level = 4'd0;
reg soc_videosoc_sdram_bankmachine0_replace = 1'd0;
reg [2:0] soc_videosoc_sdram_bankmachine0_produce = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine0_consume = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine0_wrport_adr = 3'd0;
wire [24:0] soc_videosoc_sdram_bankmachine0_wrport_dat_r;
wire soc_videosoc_sdram_bankmachine0_wrport_we;
wire [24:0] soc_videosoc_sdram_bankmachine0_wrport_dat_w;
wire soc_videosoc_sdram_bankmachine0_do_read;
wire [2:0] soc_videosoc_sdram_bankmachine0_rdport_adr;
wire [24:0] soc_videosoc_sdram_bankmachine0_rdport_dat_r;
wire soc_videosoc_sdram_bankmachine0_fifo_in_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine0_fifo_in_payload_adr;
wire soc_videosoc_sdram_bankmachine0_fifo_in_first;
wire soc_videosoc_sdram_bankmachine0_fifo_in_last;
wire soc_videosoc_sdram_bankmachine0_fifo_out_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine0_fifo_out_payload_adr;
wire soc_videosoc_sdram_bankmachine0_fifo_out_first;
wire soc_videosoc_sdram_bankmachine0_fifo_out_last;
reg soc_videosoc_sdram_bankmachine0_has_openrow = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine0_openrow = 15'd0;
wire soc_videosoc_sdram_bankmachine0_hit;
reg soc_videosoc_sdram_bankmachine0_track_open = 1'd0;
reg soc_videosoc_sdram_bankmachine0_track_close = 1'd0;
reg soc_videosoc_sdram_bankmachine0_sel_row_adr = 1'd0;
wire soc_videosoc_sdram_bankmachine0_wait;
wire soc_videosoc_sdram_bankmachine0_done;
reg [2:0] soc_videosoc_sdram_bankmachine0_count = 3'd5;
wire soc_videosoc_sdram_bankmachine1_req_valid;
wire soc_videosoc_sdram_bankmachine1_req_ready;
wire soc_videosoc_sdram_bankmachine1_req_we;
wire [21:0] soc_videosoc_sdram_bankmachine1_req_adr;
wire soc_videosoc_sdram_bankmachine1_req_lock;
reg soc_videosoc_sdram_bankmachine1_req_wdata_ready = 1'd0;
reg soc_videosoc_sdram_bankmachine1_req_rdata_valid = 1'd0;
wire soc_videosoc_sdram_bankmachine1_refresh_req;
reg soc_videosoc_sdram_bankmachine1_refresh_gnt = 1'd0;
reg soc_videosoc_sdram_bankmachine1_cmd_valid = 1'd0;
reg soc_videosoc_sdram_bankmachine1_cmd_ready = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine1_cmd_payload_a = 15'd0;
wire [2:0] soc_videosoc_sdram_bankmachine1_cmd_payload_ba;
reg soc_videosoc_sdram_bankmachine1_cmd_payload_cas = 1'd0;
reg soc_videosoc_sdram_bankmachine1_cmd_payload_ras = 1'd0;
reg soc_videosoc_sdram_bankmachine1_cmd_payload_we = 1'd0;
reg soc_videosoc_sdram_bankmachine1_cmd_payload_is_cmd = 1'd0;
reg soc_videosoc_sdram_bankmachine1_cmd_payload_is_read = 1'd0;
reg soc_videosoc_sdram_bankmachine1_cmd_payload_is_write = 1'd0;
wire soc_videosoc_sdram_bankmachine1_sink_valid;
wire soc_videosoc_sdram_bankmachine1_sink_ready;
reg soc_videosoc_sdram_bankmachine1_sink_first = 1'd0;
reg soc_videosoc_sdram_bankmachine1_sink_last = 1'd0;
wire soc_videosoc_sdram_bankmachine1_sink_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine1_sink_payload_adr;
wire soc_videosoc_sdram_bankmachine1_source_valid;
wire soc_videosoc_sdram_bankmachine1_source_ready;
wire soc_videosoc_sdram_bankmachine1_source_first;
wire soc_videosoc_sdram_bankmachine1_source_last;
wire soc_videosoc_sdram_bankmachine1_source_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine1_source_payload_adr;
wire soc_videosoc_sdram_bankmachine1_syncfifo1_we;
wire soc_videosoc_sdram_bankmachine1_syncfifo1_writable;
wire soc_videosoc_sdram_bankmachine1_syncfifo1_re;
wire soc_videosoc_sdram_bankmachine1_syncfifo1_readable;
wire [24:0] soc_videosoc_sdram_bankmachine1_syncfifo1_din;
wire [24:0] soc_videosoc_sdram_bankmachine1_syncfifo1_dout;
reg [3:0] soc_videosoc_sdram_bankmachine1_level = 4'd0;
reg soc_videosoc_sdram_bankmachine1_replace = 1'd0;
reg [2:0] soc_videosoc_sdram_bankmachine1_produce = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine1_consume = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine1_wrport_adr = 3'd0;
wire [24:0] soc_videosoc_sdram_bankmachine1_wrport_dat_r;
wire soc_videosoc_sdram_bankmachine1_wrport_we;
wire [24:0] soc_videosoc_sdram_bankmachine1_wrport_dat_w;
wire soc_videosoc_sdram_bankmachine1_do_read;
wire [2:0] soc_videosoc_sdram_bankmachine1_rdport_adr;
wire [24:0] soc_videosoc_sdram_bankmachine1_rdport_dat_r;
wire soc_videosoc_sdram_bankmachine1_fifo_in_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine1_fifo_in_payload_adr;
wire soc_videosoc_sdram_bankmachine1_fifo_in_first;
wire soc_videosoc_sdram_bankmachine1_fifo_in_last;
wire soc_videosoc_sdram_bankmachine1_fifo_out_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine1_fifo_out_payload_adr;
wire soc_videosoc_sdram_bankmachine1_fifo_out_first;
wire soc_videosoc_sdram_bankmachine1_fifo_out_last;
reg soc_videosoc_sdram_bankmachine1_has_openrow = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine1_openrow = 15'd0;
wire soc_videosoc_sdram_bankmachine1_hit;
reg soc_videosoc_sdram_bankmachine1_track_open = 1'd0;
reg soc_videosoc_sdram_bankmachine1_track_close = 1'd0;
reg soc_videosoc_sdram_bankmachine1_sel_row_adr = 1'd0;
wire soc_videosoc_sdram_bankmachine1_wait;
wire soc_videosoc_sdram_bankmachine1_done;
reg [2:0] soc_videosoc_sdram_bankmachine1_count = 3'd5;
wire soc_videosoc_sdram_bankmachine2_req_valid;
wire soc_videosoc_sdram_bankmachine2_req_ready;
wire soc_videosoc_sdram_bankmachine2_req_we;
wire [21:0] soc_videosoc_sdram_bankmachine2_req_adr;
wire soc_videosoc_sdram_bankmachine2_req_lock;
reg soc_videosoc_sdram_bankmachine2_req_wdata_ready = 1'd0;
reg soc_videosoc_sdram_bankmachine2_req_rdata_valid = 1'd0;
wire soc_videosoc_sdram_bankmachine2_refresh_req;
reg soc_videosoc_sdram_bankmachine2_refresh_gnt = 1'd0;
reg soc_videosoc_sdram_bankmachine2_cmd_valid = 1'd0;
reg soc_videosoc_sdram_bankmachine2_cmd_ready = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine2_cmd_payload_a = 15'd0;
wire [2:0] soc_videosoc_sdram_bankmachine2_cmd_payload_ba;
reg soc_videosoc_sdram_bankmachine2_cmd_payload_cas = 1'd0;
reg soc_videosoc_sdram_bankmachine2_cmd_payload_ras = 1'd0;
reg soc_videosoc_sdram_bankmachine2_cmd_payload_we = 1'd0;
reg soc_videosoc_sdram_bankmachine2_cmd_payload_is_cmd = 1'd0;
reg soc_videosoc_sdram_bankmachine2_cmd_payload_is_read = 1'd0;
reg soc_videosoc_sdram_bankmachine2_cmd_payload_is_write = 1'd0;
wire soc_videosoc_sdram_bankmachine2_sink_valid;
wire soc_videosoc_sdram_bankmachine2_sink_ready;
reg soc_videosoc_sdram_bankmachine2_sink_first = 1'd0;
reg soc_videosoc_sdram_bankmachine2_sink_last = 1'd0;
wire soc_videosoc_sdram_bankmachine2_sink_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine2_sink_payload_adr;
wire soc_videosoc_sdram_bankmachine2_source_valid;
wire soc_videosoc_sdram_bankmachine2_source_ready;
wire soc_videosoc_sdram_bankmachine2_source_first;
wire soc_videosoc_sdram_bankmachine2_source_last;
wire soc_videosoc_sdram_bankmachine2_source_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine2_source_payload_adr;
wire soc_videosoc_sdram_bankmachine2_syncfifo2_we;
wire soc_videosoc_sdram_bankmachine2_syncfifo2_writable;
wire soc_videosoc_sdram_bankmachine2_syncfifo2_re;
wire soc_videosoc_sdram_bankmachine2_syncfifo2_readable;
wire [24:0] soc_videosoc_sdram_bankmachine2_syncfifo2_din;
wire [24:0] soc_videosoc_sdram_bankmachine2_syncfifo2_dout;
reg [3:0] soc_videosoc_sdram_bankmachine2_level = 4'd0;
reg soc_videosoc_sdram_bankmachine2_replace = 1'd0;
reg [2:0] soc_videosoc_sdram_bankmachine2_produce = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine2_consume = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine2_wrport_adr = 3'd0;
wire [24:0] soc_videosoc_sdram_bankmachine2_wrport_dat_r;
wire soc_videosoc_sdram_bankmachine2_wrport_we;
wire [24:0] soc_videosoc_sdram_bankmachine2_wrport_dat_w;
wire soc_videosoc_sdram_bankmachine2_do_read;
wire [2:0] soc_videosoc_sdram_bankmachine2_rdport_adr;
wire [24:0] soc_videosoc_sdram_bankmachine2_rdport_dat_r;
wire soc_videosoc_sdram_bankmachine2_fifo_in_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine2_fifo_in_payload_adr;
wire soc_videosoc_sdram_bankmachine2_fifo_in_first;
wire soc_videosoc_sdram_bankmachine2_fifo_in_last;
wire soc_videosoc_sdram_bankmachine2_fifo_out_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine2_fifo_out_payload_adr;
wire soc_videosoc_sdram_bankmachine2_fifo_out_first;
wire soc_videosoc_sdram_bankmachine2_fifo_out_last;
reg soc_videosoc_sdram_bankmachine2_has_openrow = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine2_openrow = 15'd0;
wire soc_videosoc_sdram_bankmachine2_hit;
reg soc_videosoc_sdram_bankmachine2_track_open = 1'd0;
reg soc_videosoc_sdram_bankmachine2_track_close = 1'd0;
reg soc_videosoc_sdram_bankmachine2_sel_row_adr = 1'd0;
wire soc_videosoc_sdram_bankmachine2_wait;
wire soc_videosoc_sdram_bankmachine2_done;
reg [2:0] soc_videosoc_sdram_bankmachine2_count = 3'd5;
wire soc_videosoc_sdram_bankmachine3_req_valid;
wire soc_videosoc_sdram_bankmachine3_req_ready;
wire soc_videosoc_sdram_bankmachine3_req_we;
wire [21:0] soc_videosoc_sdram_bankmachine3_req_adr;
wire soc_videosoc_sdram_bankmachine3_req_lock;
reg soc_videosoc_sdram_bankmachine3_req_wdata_ready = 1'd0;
reg soc_videosoc_sdram_bankmachine3_req_rdata_valid = 1'd0;
wire soc_videosoc_sdram_bankmachine3_refresh_req;
reg soc_videosoc_sdram_bankmachine3_refresh_gnt = 1'd0;
reg soc_videosoc_sdram_bankmachine3_cmd_valid = 1'd0;
reg soc_videosoc_sdram_bankmachine3_cmd_ready = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine3_cmd_payload_a = 15'd0;
wire [2:0] soc_videosoc_sdram_bankmachine3_cmd_payload_ba;
reg soc_videosoc_sdram_bankmachine3_cmd_payload_cas = 1'd0;
reg soc_videosoc_sdram_bankmachine3_cmd_payload_ras = 1'd0;
reg soc_videosoc_sdram_bankmachine3_cmd_payload_we = 1'd0;
reg soc_videosoc_sdram_bankmachine3_cmd_payload_is_cmd = 1'd0;
reg soc_videosoc_sdram_bankmachine3_cmd_payload_is_read = 1'd0;
reg soc_videosoc_sdram_bankmachine3_cmd_payload_is_write = 1'd0;
wire soc_videosoc_sdram_bankmachine3_sink_valid;
wire soc_videosoc_sdram_bankmachine3_sink_ready;
reg soc_videosoc_sdram_bankmachine3_sink_first = 1'd0;
reg soc_videosoc_sdram_bankmachine3_sink_last = 1'd0;
wire soc_videosoc_sdram_bankmachine3_sink_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine3_sink_payload_adr;
wire soc_videosoc_sdram_bankmachine3_source_valid;
wire soc_videosoc_sdram_bankmachine3_source_ready;
wire soc_videosoc_sdram_bankmachine3_source_first;
wire soc_videosoc_sdram_bankmachine3_source_last;
wire soc_videosoc_sdram_bankmachine3_source_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine3_source_payload_adr;
wire soc_videosoc_sdram_bankmachine3_syncfifo3_we;
wire soc_videosoc_sdram_bankmachine3_syncfifo3_writable;
wire soc_videosoc_sdram_bankmachine3_syncfifo3_re;
wire soc_videosoc_sdram_bankmachine3_syncfifo3_readable;
wire [24:0] soc_videosoc_sdram_bankmachine3_syncfifo3_din;
wire [24:0] soc_videosoc_sdram_bankmachine3_syncfifo3_dout;
reg [3:0] soc_videosoc_sdram_bankmachine3_level = 4'd0;
reg soc_videosoc_sdram_bankmachine3_replace = 1'd0;
reg [2:0] soc_videosoc_sdram_bankmachine3_produce = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine3_consume = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine3_wrport_adr = 3'd0;
wire [24:0] soc_videosoc_sdram_bankmachine3_wrport_dat_r;
wire soc_videosoc_sdram_bankmachine3_wrport_we;
wire [24:0] soc_videosoc_sdram_bankmachine3_wrport_dat_w;
wire soc_videosoc_sdram_bankmachine3_do_read;
wire [2:0] soc_videosoc_sdram_bankmachine3_rdport_adr;
wire [24:0] soc_videosoc_sdram_bankmachine3_rdport_dat_r;
wire soc_videosoc_sdram_bankmachine3_fifo_in_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine3_fifo_in_payload_adr;
wire soc_videosoc_sdram_bankmachine3_fifo_in_first;
wire soc_videosoc_sdram_bankmachine3_fifo_in_last;
wire soc_videosoc_sdram_bankmachine3_fifo_out_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine3_fifo_out_payload_adr;
wire soc_videosoc_sdram_bankmachine3_fifo_out_first;
wire soc_videosoc_sdram_bankmachine3_fifo_out_last;
reg soc_videosoc_sdram_bankmachine3_has_openrow = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine3_openrow = 15'd0;
wire soc_videosoc_sdram_bankmachine3_hit;
reg soc_videosoc_sdram_bankmachine3_track_open = 1'd0;
reg soc_videosoc_sdram_bankmachine3_track_close = 1'd0;
reg soc_videosoc_sdram_bankmachine3_sel_row_adr = 1'd0;
wire soc_videosoc_sdram_bankmachine3_wait;
wire soc_videosoc_sdram_bankmachine3_done;
reg [2:0] soc_videosoc_sdram_bankmachine3_count = 3'd5;
wire soc_videosoc_sdram_bankmachine4_req_valid;
wire soc_videosoc_sdram_bankmachine4_req_ready;
wire soc_videosoc_sdram_bankmachine4_req_we;
wire [21:0] soc_videosoc_sdram_bankmachine4_req_adr;
wire soc_videosoc_sdram_bankmachine4_req_lock;
reg soc_videosoc_sdram_bankmachine4_req_wdata_ready = 1'd0;
reg soc_videosoc_sdram_bankmachine4_req_rdata_valid = 1'd0;
wire soc_videosoc_sdram_bankmachine4_refresh_req;
reg soc_videosoc_sdram_bankmachine4_refresh_gnt = 1'd0;
reg soc_videosoc_sdram_bankmachine4_cmd_valid = 1'd0;
reg soc_videosoc_sdram_bankmachine4_cmd_ready = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine4_cmd_payload_a = 15'd0;
wire [2:0] soc_videosoc_sdram_bankmachine4_cmd_payload_ba;
reg soc_videosoc_sdram_bankmachine4_cmd_payload_cas = 1'd0;
reg soc_videosoc_sdram_bankmachine4_cmd_payload_ras = 1'd0;
reg soc_videosoc_sdram_bankmachine4_cmd_payload_we = 1'd0;
reg soc_videosoc_sdram_bankmachine4_cmd_payload_is_cmd = 1'd0;
reg soc_videosoc_sdram_bankmachine4_cmd_payload_is_read = 1'd0;
reg soc_videosoc_sdram_bankmachine4_cmd_payload_is_write = 1'd0;
wire soc_videosoc_sdram_bankmachine4_sink_valid;
wire soc_videosoc_sdram_bankmachine4_sink_ready;
reg soc_videosoc_sdram_bankmachine4_sink_first = 1'd0;
reg soc_videosoc_sdram_bankmachine4_sink_last = 1'd0;
wire soc_videosoc_sdram_bankmachine4_sink_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine4_sink_payload_adr;
wire soc_videosoc_sdram_bankmachine4_source_valid;
wire soc_videosoc_sdram_bankmachine4_source_ready;
wire soc_videosoc_sdram_bankmachine4_source_first;
wire soc_videosoc_sdram_bankmachine4_source_last;
wire soc_videosoc_sdram_bankmachine4_source_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine4_source_payload_adr;
wire soc_videosoc_sdram_bankmachine4_syncfifo4_we;
wire soc_videosoc_sdram_bankmachine4_syncfifo4_writable;
wire soc_videosoc_sdram_bankmachine4_syncfifo4_re;
wire soc_videosoc_sdram_bankmachine4_syncfifo4_readable;
wire [24:0] soc_videosoc_sdram_bankmachine4_syncfifo4_din;
wire [24:0] soc_videosoc_sdram_bankmachine4_syncfifo4_dout;
reg [3:0] soc_videosoc_sdram_bankmachine4_level = 4'd0;
reg soc_videosoc_sdram_bankmachine4_replace = 1'd0;
reg [2:0] soc_videosoc_sdram_bankmachine4_produce = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine4_consume = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine4_wrport_adr = 3'd0;
wire [24:0] soc_videosoc_sdram_bankmachine4_wrport_dat_r;
wire soc_videosoc_sdram_bankmachine4_wrport_we;
wire [24:0] soc_videosoc_sdram_bankmachine4_wrport_dat_w;
wire soc_videosoc_sdram_bankmachine4_do_read;
wire [2:0] soc_videosoc_sdram_bankmachine4_rdport_adr;
wire [24:0] soc_videosoc_sdram_bankmachine4_rdport_dat_r;
wire soc_videosoc_sdram_bankmachine4_fifo_in_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine4_fifo_in_payload_adr;
wire soc_videosoc_sdram_bankmachine4_fifo_in_first;
wire soc_videosoc_sdram_bankmachine4_fifo_in_last;
wire soc_videosoc_sdram_bankmachine4_fifo_out_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine4_fifo_out_payload_adr;
wire soc_videosoc_sdram_bankmachine4_fifo_out_first;
wire soc_videosoc_sdram_bankmachine4_fifo_out_last;
reg soc_videosoc_sdram_bankmachine4_has_openrow = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine4_openrow = 15'd0;
wire soc_videosoc_sdram_bankmachine4_hit;
reg soc_videosoc_sdram_bankmachine4_track_open = 1'd0;
reg soc_videosoc_sdram_bankmachine4_track_close = 1'd0;
reg soc_videosoc_sdram_bankmachine4_sel_row_adr = 1'd0;
wire soc_videosoc_sdram_bankmachine4_wait;
wire soc_videosoc_sdram_bankmachine4_done;
reg [2:0] soc_videosoc_sdram_bankmachine4_count = 3'd5;
wire soc_videosoc_sdram_bankmachine5_req_valid;
wire soc_videosoc_sdram_bankmachine5_req_ready;
wire soc_videosoc_sdram_bankmachine5_req_we;
wire [21:0] soc_videosoc_sdram_bankmachine5_req_adr;
wire soc_videosoc_sdram_bankmachine5_req_lock;
reg soc_videosoc_sdram_bankmachine5_req_wdata_ready = 1'd0;
reg soc_videosoc_sdram_bankmachine5_req_rdata_valid = 1'd0;
wire soc_videosoc_sdram_bankmachine5_refresh_req;
reg soc_videosoc_sdram_bankmachine5_refresh_gnt = 1'd0;
reg soc_videosoc_sdram_bankmachine5_cmd_valid = 1'd0;
reg soc_videosoc_sdram_bankmachine5_cmd_ready = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine5_cmd_payload_a = 15'd0;
wire [2:0] soc_videosoc_sdram_bankmachine5_cmd_payload_ba;
reg soc_videosoc_sdram_bankmachine5_cmd_payload_cas = 1'd0;
reg soc_videosoc_sdram_bankmachine5_cmd_payload_ras = 1'd0;
reg soc_videosoc_sdram_bankmachine5_cmd_payload_we = 1'd0;
reg soc_videosoc_sdram_bankmachine5_cmd_payload_is_cmd = 1'd0;
reg soc_videosoc_sdram_bankmachine5_cmd_payload_is_read = 1'd0;
reg soc_videosoc_sdram_bankmachine5_cmd_payload_is_write = 1'd0;
wire soc_videosoc_sdram_bankmachine5_sink_valid;
wire soc_videosoc_sdram_bankmachine5_sink_ready;
reg soc_videosoc_sdram_bankmachine5_sink_first = 1'd0;
reg soc_videosoc_sdram_bankmachine5_sink_last = 1'd0;
wire soc_videosoc_sdram_bankmachine5_sink_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine5_sink_payload_adr;
wire soc_videosoc_sdram_bankmachine5_source_valid;
wire soc_videosoc_sdram_bankmachine5_source_ready;
wire soc_videosoc_sdram_bankmachine5_source_first;
wire soc_videosoc_sdram_bankmachine5_source_last;
wire soc_videosoc_sdram_bankmachine5_source_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine5_source_payload_adr;
wire soc_videosoc_sdram_bankmachine5_syncfifo5_we;
wire soc_videosoc_sdram_bankmachine5_syncfifo5_writable;
wire soc_videosoc_sdram_bankmachine5_syncfifo5_re;
wire soc_videosoc_sdram_bankmachine5_syncfifo5_readable;
wire [24:0] soc_videosoc_sdram_bankmachine5_syncfifo5_din;
wire [24:0] soc_videosoc_sdram_bankmachine5_syncfifo5_dout;
reg [3:0] soc_videosoc_sdram_bankmachine5_level = 4'd0;
reg soc_videosoc_sdram_bankmachine5_replace = 1'd0;
reg [2:0] soc_videosoc_sdram_bankmachine5_produce = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine5_consume = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine5_wrport_adr = 3'd0;
wire [24:0] soc_videosoc_sdram_bankmachine5_wrport_dat_r;
wire soc_videosoc_sdram_bankmachine5_wrport_we;
wire [24:0] soc_videosoc_sdram_bankmachine5_wrport_dat_w;
wire soc_videosoc_sdram_bankmachine5_do_read;
wire [2:0] soc_videosoc_sdram_bankmachine5_rdport_adr;
wire [24:0] soc_videosoc_sdram_bankmachine5_rdport_dat_r;
wire soc_videosoc_sdram_bankmachine5_fifo_in_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine5_fifo_in_payload_adr;
wire soc_videosoc_sdram_bankmachine5_fifo_in_first;
wire soc_videosoc_sdram_bankmachine5_fifo_in_last;
wire soc_videosoc_sdram_bankmachine5_fifo_out_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine5_fifo_out_payload_adr;
wire soc_videosoc_sdram_bankmachine5_fifo_out_first;
wire soc_videosoc_sdram_bankmachine5_fifo_out_last;
reg soc_videosoc_sdram_bankmachine5_has_openrow = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine5_openrow = 15'd0;
wire soc_videosoc_sdram_bankmachine5_hit;
reg soc_videosoc_sdram_bankmachine5_track_open = 1'd0;
reg soc_videosoc_sdram_bankmachine5_track_close = 1'd0;
reg soc_videosoc_sdram_bankmachine5_sel_row_adr = 1'd0;
wire soc_videosoc_sdram_bankmachine5_wait;
wire soc_videosoc_sdram_bankmachine5_done;
reg [2:0] soc_videosoc_sdram_bankmachine5_count = 3'd5;
wire soc_videosoc_sdram_bankmachine6_req_valid;
wire soc_videosoc_sdram_bankmachine6_req_ready;
wire soc_videosoc_sdram_bankmachine6_req_we;
wire [21:0] soc_videosoc_sdram_bankmachine6_req_adr;
wire soc_videosoc_sdram_bankmachine6_req_lock;
reg soc_videosoc_sdram_bankmachine6_req_wdata_ready = 1'd0;
reg soc_videosoc_sdram_bankmachine6_req_rdata_valid = 1'd0;
wire soc_videosoc_sdram_bankmachine6_refresh_req;
reg soc_videosoc_sdram_bankmachine6_refresh_gnt = 1'd0;
reg soc_videosoc_sdram_bankmachine6_cmd_valid = 1'd0;
reg soc_videosoc_sdram_bankmachine6_cmd_ready = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine6_cmd_payload_a = 15'd0;
wire [2:0] soc_videosoc_sdram_bankmachine6_cmd_payload_ba;
reg soc_videosoc_sdram_bankmachine6_cmd_payload_cas = 1'd0;
reg soc_videosoc_sdram_bankmachine6_cmd_payload_ras = 1'd0;
reg soc_videosoc_sdram_bankmachine6_cmd_payload_we = 1'd0;
reg soc_videosoc_sdram_bankmachine6_cmd_payload_is_cmd = 1'd0;
reg soc_videosoc_sdram_bankmachine6_cmd_payload_is_read = 1'd0;
reg soc_videosoc_sdram_bankmachine6_cmd_payload_is_write = 1'd0;
wire soc_videosoc_sdram_bankmachine6_sink_valid;
wire soc_videosoc_sdram_bankmachine6_sink_ready;
reg soc_videosoc_sdram_bankmachine6_sink_first = 1'd0;
reg soc_videosoc_sdram_bankmachine6_sink_last = 1'd0;
wire soc_videosoc_sdram_bankmachine6_sink_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine6_sink_payload_adr;
wire soc_videosoc_sdram_bankmachine6_source_valid;
wire soc_videosoc_sdram_bankmachine6_source_ready;
wire soc_videosoc_sdram_bankmachine6_source_first;
wire soc_videosoc_sdram_bankmachine6_source_last;
wire soc_videosoc_sdram_bankmachine6_source_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine6_source_payload_adr;
wire soc_videosoc_sdram_bankmachine6_syncfifo6_we;
wire soc_videosoc_sdram_bankmachine6_syncfifo6_writable;
wire soc_videosoc_sdram_bankmachine6_syncfifo6_re;
wire soc_videosoc_sdram_bankmachine6_syncfifo6_readable;
wire [24:0] soc_videosoc_sdram_bankmachine6_syncfifo6_din;
wire [24:0] soc_videosoc_sdram_bankmachine6_syncfifo6_dout;
reg [3:0] soc_videosoc_sdram_bankmachine6_level = 4'd0;
reg soc_videosoc_sdram_bankmachine6_replace = 1'd0;
reg [2:0] soc_videosoc_sdram_bankmachine6_produce = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine6_consume = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine6_wrport_adr = 3'd0;
wire [24:0] soc_videosoc_sdram_bankmachine6_wrport_dat_r;
wire soc_videosoc_sdram_bankmachine6_wrport_we;
wire [24:0] soc_videosoc_sdram_bankmachine6_wrport_dat_w;
wire soc_videosoc_sdram_bankmachine6_do_read;
wire [2:0] soc_videosoc_sdram_bankmachine6_rdport_adr;
wire [24:0] soc_videosoc_sdram_bankmachine6_rdport_dat_r;
wire soc_videosoc_sdram_bankmachine6_fifo_in_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine6_fifo_in_payload_adr;
wire soc_videosoc_sdram_bankmachine6_fifo_in_first;
wire soc_videosoc_sdram_bankmachine6_fifo_in_last;
wire soc_videosoc_sdram_bankmachine6_fifo_out_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine6_fifo_out_payload_adr;
wire soc_videosoc_sdram_bankmachine6_fifo_out_first;
wire soc_videosoc_sdram_bankmachine6_fifo_out_last;
reg soc_videosoc_sdram_bankmachine6_has_openrow = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine6_openrow = 15'd0;
wire soc_videosoc_sdram_bankmachine6_hit;
reg soc_videosoc_sdram_bankmachine6_track_open = 1'd0;
reg soc_videosoc_sdram_bankmachine6_track_close = 1'd0;
reg soc_videosoc_sdram_bankmachine6_sel_row_adr = 1'd0;
wire soc_videosoc_sdram_bankmachine6_wait;
wire soc_videosoc_sdram_bankmachine6_done;
reg [2:0] soc_videosoc_sdram_bankmachine6_count = 3'd5;
wire soc_videosoc_sdram_bankmachine7_req_valid;
wire soc_videosoc_sdram_bankmachine7_req_ready;
wire soc_videosoc_sdram_bankmachine7_req_we;
wire [21:0] soc_videosoc_sdram_bankmachine7_req_adr;
wire soc_videosoc_sdram_bankmachine7_req_lock;
reg soc_videosoc_sdram_bankmachine7_req_wdata_ready = 1'd0;
reg soc_videosoc_sdram_bankmachine7_req_rdata_valid = 1'd0;
wire soc_videosoc_sdram_bankmachine7_refresh_req;
reg soc_videosoc_sdram_bankmachine7_refresh_gnt = 1'd0;
reg soc_videosoc_sdram_bankmachine7_cmd_valid = 1'd0;
reg soc_videosoc_sdram_bankmachine7_cmd_ready = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine7_cmd_payload_a = 15'd0;
wire [2:0] soc_videosoc_sdram_bankmachine7_cmd_payload_ba;
reg soc_videosoc_sdram_bankmachine7_cmd_payload_cas = 1'd0;
reg soc_videosoc_sdram_bankmachine7_cmd_payload_ras = 1'd0;
reg soc_videosoc_sdram_bankmachine7_cmd_payload_we = 1'd0;
reg soc_videosoc_sdram_bankmachine7_cmd_payload_is_cmd = 1'd0;
reg soc_videosoc_sdram_bankmachine7_cmd_payload_is_read = 1'd0;
reg soc_videosoc_sdram_bankmachine7_cmd_payload_is_write = 1'd0;
wire soc_videosoc_sdram_bankmachine7_sink_valid;
wire soc_videosoc_sdram_bankmachine7_sink_ready;
reg soc_videosoc_sdram_bankmachine7_sink_first = 1'd0;
reg soc_videosoc_sdram_bankmachine7_sink_last = 1'd0;
wire soc_videosoc_sdram_bankmachine7_sink_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine7_sink_payload_adr;
wire soc_videosoc_sdram_bankmachine7_source_valid;
wire soc_videosoc_sdram_bankmachine7_source_ready;
wire soc_videosoc_sdram_bankmachine7_source_first;
wire soc_videosoc_sdram_bankmachine7_source_last;
wire soc_videosoc_sdram_bankmachine7_source_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine7_source_payload_adr;
wire soc_videosoc_sdram_bankmachine7_syncfifo7_we;
wire soc_videosoc_sdram_bankmachine7_syncfifo7_writable;
wire soc_videosoc_sdram_bankmachine7_syncfifo7_re;
wire soc_videosoc_sdram_bankmachine7_syncfifo7_readable;
wire [24:0] soc_videosoc_sdram_bankmachine7_syncfifo7_din;
wire [24:0] soc_videosoc_sdram_bankmachine7_syncfifo7_dout;
reg [3:0] soc_videosoc_sdram_bankmachine7_level = 4'd0;
reg soc_videosoc_sdram_bankmachine7_replace = 1'd0;
reg [2:0] soc_videosoc_sdram_bankmachine7_produce = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine7_consume = 3'd0;
reg [2:0] soc_videosoc_sdram_bankmachine7_wrport_adr = 3'd0;
wire [24:0] soc_videosoc_sdram_bankmachine7_wrport_dat_r;
wire soc_videosoc_sdram_bankmachine7_wrport_we;
wire [24:0] soc_videosoc_sdram_bankmachine7_wrport_dat_w;
wire soc_videosoc_sdram_bankmachine7_do_read;
wire [2:0] soc_videosoc_sdram_bankmachine7_rdport_adr;
wire [24:0] soc_videosoc_sdram_bankmachine7_rdport_dat_r;
wire soc_videosoc_sdram_bankmachine7_fifo_in_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine7_fifo_in_payload_adr;
wire soc_videosoc_sdram_bankmachine7_fifo_in_first;
wire soc_videosoc_sdram_bankmachine7_fifo_in_last;
wire soc_videosoc_sdram_bankmachine7_fifo_out_payload_we;
wire [21:0] soc_videosoc_sdram_bankmachine7_fifo_out_payload_adr;
wire soc_videosoc_sdram_bankmachine7_fifo_out_first;
wire soc_videosoc_sdram_bankmachine7_fifo_out_last;
reg soc_videosoc_sdram_bankmachine7_has_openrow = 1'd0;
reg [14:0] soc_videosoc_sdram_bankmachine7_openrow = 15'd0;
wire soc_videosoc_sdram_bankmachine7_hit;
reg soc_videosoc_sdram_bankmachine7_track_open = 1'd0;
reg soc_videosoc_sdram_bankmachine7_track_close = 1'd0;
reg soc_videosoc_sdram_bankmachine7_sel_row_adr = 1'd0;
wire soc_videosoc_sdram_bankmachine7_wait;
wire soc_videosoc_sdram_bankmachine7_done;
reg [2:0] soc_videosoc_sdram_bankmachine7_count = 3'd5;
reg soc_videosoc_sdram_choose_cmd_want_reads = 1'd0;
reg soc_videosoc_sdram_choose_cmd_want_writes = 1'd0;
reg soc_videosoc_sdram_choose_cmd_want_cmds = 1'd0;
wire soc_videosoc_sdram_choose_cmd_cmd_valid;
reg soc_videosoc_sdram_choose_cmd_cmd_ready = 1'd0;
wire [14:0] soc_videosoc_sdram_choose_cmd_cmd_payload_a;
wire [2:0] soc_videosoc_sdram_choose_cmd_cmd_payload_ba;
reg soc_videosoc_sdram_choose_cmd_cmd_payload_cas = 1'd0;
reg soc_videosoc_sdram_choose_cmd_cmd_payload_ras = 1'd0;
reg soc_videosoc_sdram_choose_cmd_cmd_payload_we = 1'd0;
wire soc_videosoc_sdram_choose_cmd_cmd_payload_is_cmd;
wire soc_videosoc_sdram_choose_cmd_cmd_payload_is_read;
wire soc_videosoc_sdram_choose_cmd_cmd_payload_is_write;
reg [7:0] soc_videosoc_sdram_choose_cmd_valids = 8'd0;
wire [7:0] soc_videosoc_sdram_choose_cmd_request;
reg [2:0] soc_videosoc_sdram_choose_cmd_grant = 3'd0;
wire soc_videosoc_sdram_choose_cmd_ce;
reg soc_videosoc_sdram_choose_req_want_reads = 1'd0;
reg soc_videosoc_sdram_choose_req_want_writes = 1'd0;
reg soc_videosoc_sdram_choose_req_want_cmds = 1'd0;
wire soc_videosoc_sdram_choose_req_cmd_valid;
reg soc_videosoc_sdram_choose_req_cmd_ready = 1'd0;
wire [14:0] soc_videosoc_sdram_choose_req_cmd_payload_a;
wire [2:0] soc_videosoc_sdram_choose_req_cmd_payload_ba;
reg soc_videosoc_sdram_choose_req_cmd_payload_cas = 1'd0;
reg soc_videosoc_sdram_choose_req_cmd_payload_ras = 1'd0;
reg soc_videosoc_sdram_choose_req_cmd_payload_we = 1'd0;
wire soc_videosoc_sdram_choose_req_cmd_payload_is_cmd;
wire soc_videosoc_sdram_choose_req_cmd_payload_is_read;
wire soc_videosoc_sdram_choose_req_cmd_payload_is_write;
reg [7:0] soc_videosoc_sdram_choose_req_valids = 8'd0;
wire [7:0] soc_videosoc_sdram_choose_req_request;
reg [2:0] soc_videosoc_sdram_choose_req_grant = 3'd0;
wire soc_videosoc_sdram_choose_req_ce;
reg [14:0] soc_videosoc_sdram_nop_a = 15'd0;
reg [2:0] soc_videosoc_sdram_nop_ba = 3'd0;
reg soc_videosoc_sdram_nop_cas = 1'd0;
reg soc_videosoc_sdram_nop_ras = 1'd0;
reg soc_videosoc_sdram_nop_we = 1'd0;
reg [1:0] soc_videosoc_sdram_sel0 = 2'd0;
reg [1:0] soc_videosoc_sdram_sel1 = 2'd0;
reg [1:0] soc_videosoc_sdram_sel2 = 2'd0;
reg [1:0] soc_videosoc_sdram_sel3 = 2'd0;
wire soc_videosoc_sdram_read_available;
wire soc_videosoc_sdram_write_available;
reg soc_videosoc_sdram_en0 = 1'd0;
wire soc_videosoc_sdram_max_time0;
reg [4:0] soc_videosoc_sdram_time0 = 5'd0;
reg soc_videosoc_sdram_en1 = 1'd0;
wire soc_videosoc_sdram_max_time1;
reg [3:0] soc_videosoc_sdram_time1 = 4'd0;
wire soc_videosoc_sdram_go_to_refresh;
wire soc_videosoc_sdram_bandwidth_update_re;
wire soc_videosoc_sdram_bandwidth_update_r;
reg soc_videosoc_sdram_bandwidth_update_w = 1'd0;
reg [23:0] soc_videosoc_sdram_bandwidth_nreads_status = 24'd0;
reg [23:0] soc_videosoc_sdram_bandwidth_nwrites_status = 24'd0;
reg [7:0] soc_videosoc_sdram_bandwidth_data_width_status = 8'd128;
reg soc_videosoc_sdram_bandwidth_cmd_valid = 1'd0;
reg soc_videosoc_sdram_bandwidth_cmd_ready = 1'd0;
reg soc_videosoc_sdram_bandwidth_cmd_is_read = 1'd0;
reg soc_videosoc_sdram_bandwidth_cmd_is_write = 1'd0;
reg [23:0] soc_videosoc_sdram_bandwidth_counter = 24'd0;
reg soc_videosoc_sdram_bandwidth_period = 1'd0;
reg [23:0] soc_videosoc_sdram_bandwidth_nreads = 24'd0;
reg [23:0] soc_videosoc_sdram_bandwidth_nwrites = 24'd0;
reg [23:0] soc_videosoc_sdram_bandwidth_nreads_r = 24'd0;
reg [23:0] soc_videosoc_sdram_bandwidth_nwrites_r = 24'd0;
wire [29:0] soc_videosoc_interface1_wb_sdram_adr;
wire [31:0] soc_videosoc_interface1_wb_sdram_dat_w;
wire [31:0] soc_videosoc_interface1_wb_sdram_dat_r;
wire [3:0] soc_videosoc_interface1_wb_sdram_sel;
wire soc_videosoc_interface1_wb_sdram_cyc;
wire soc_videosoc_interface1_wb_sdram_stb;
wire soc_videosoc_interface1_wb_sdram_ack;
wire soc_videosoc_interface1_wb_sdram_we;
wire [2:0] soc_videosoc_interface1_wb_sdram_cti;
wire [1:0] soc_videosoc_interface1_wb_sdram_bte;
wire soc_videosoc_interface1_wb_sdram_err;
reg soc_videosoc_port_cmd_valid = 1'd0;
wire soc_videosoc_port_cmd_ready;
reg soc_videosoc_port_cmd_payload_we = 1'd0;
wire [24:0] soc_videosoc_port_cmd_payload_adr;
reg soc_videosoc_port_wdata_valid = 1'd0;
wire soc_videosoc_port_wdata_ready;
wire [127:0] soc_videosoc_port_wdata_payload_data;
wire [15:0] soc_videosoc_port_wdata_payload_we;
wire soc_videosoc_port_rdata_valid;
reg soc_videosoc_port_rdata_ready = 1'd0;
wire [127:0] soc_videosoc_port_rdata_payload_data;
wire [29:0] soc_videosoc_interface_adr;
wire [127:0] soc_videosoc_interface_dat_w;
wire [127:0] soc_videosoc_interface_dat_r;
wire [15:0] soc_videosoc_interface_sel;
reg soc_videosoc_interface_cyc = 1'd0;
reg soc_videosoc_interface_stb = 1'd0;
reg soc_videosoc_interface_ack = 1'd0;
reg soc_videosoc_interface_we = 1'd0;
wire [8:0] soc_videosoc_data_port_adr;
wire [127:0] soc_videosoc_data_port_dat_r;
reg [15:0] soc_videosoc_data_port_we = 16'd0;
reg [127:0] soc_videosoc_data_port_dat_w = 128'd0;
reg soc_videosoc_write_from_slave = 1'd0;
reg [1:0] soc_videosoc_adr_offset_r = 2'd0;
wire [8:0] soc_videosoc_tag_port_adr;
wire [23:0] soc_videosoc_tag_port_dat_r;
reg soc_videosoc_tag_port_we = 1'd0;
wire [23:0] soc_videosoc_tag_port_dat_w;
wire [22:0] soc_videosoc_tag_do_tag;
wire soc_videosoc_tag_do_dirty;
wire [22:0] soc_videosoc_tag_di_tag;
reg soc_videosoc_tag_di_dirty = 1'd0;
reg soc_videosoc_word_clr = 1'd0;
reg soc_videosoc_word_inc = 1'd0;
reg soc_videosoc_clk0 = 1'd0;
wire [29:0] soc_videosoc_bus_adr;
wire [31:0] soc_videosoc_bus_dat_w;
wire [31:0] soc_videosoc_bus_dat_r;
wire [3:0] soc_videosoc_bus_sel;
wire soc_videosoc_bus_cyc;
wire soc_videosoc_bus_stb;
reg soc_videosoc_bus_ack = 1'd0;
wire soc_videosoc_bus_we;
wire [2:0] soc_videosoc_bus_cti;
wire [1:0] soc_videosoc_bus_bte;
reg soc_videosoc_bus_err = 1'd0;
reg [3:0] soc_videosoc_bitbang_storage_full = 4'd0;
wire [3:0] soc_videosoc_bitbang_storage;
reg soc_videosoc_bitbang_re = 1'd0;
reg soc_videosoc_miso_status = 1'd0;
reg soc_videosoc_bitbang_en_storage_full = 1'd0;
wire soc_videosoc_bitbang_en_storage;
reg soc_videosoc_bitbang_en_re = 1'd0;
reg soc_videosoc_cs_n = 1'd1;
reg soc_videosoc_clk1 = 1'd0;
reg [31:0] soc_videosoc_sr = 32'd0;
reg soc_videosoc_i = 1'd0;
reg soc_videosoc_miso = 1'd0;
reg [7:0] soc_videosoc_counter = 8'd0;
reg soc_ethphy_reset_storage_full = 1'd0;
wire soc_ethphy_reset_storage;
reg soc_ethphy_reset_re = 1'd0;
(* dont_touch = "true" *) wire eth_rx_clk;
wire eth_rx_rst;
(* dont_touch = "true" *) wire eth_tx_clk;
wire eth_tx_rst;
wire eth_tx90_clk;
wire soc_ethphy_eth_rx_clk_ibuf;
wire soc_ethphy_pll_locked;
wire soc_ethphy_pll_fb;
wire soc_ethphy_pll_clk_tx;
wire soc_ethphy_pll_clk_tx90;
wire soc_ethphy_eth_tx_clk_obuf;
(* ars_false_path = "true" *) wire soc_ethphy_reset0;
wire soc_ethphy_reset1;
reg [8:0] soc_ethphy_counter = 9'd0;
wire soc_ethphy_counter_done;
wire soc_ethphy_counter_ce;
wire soc_ethphy_sink_valid;
wire soc_ethphy_sink_ready;
wire soc_ethphy_sink_first;
wire soc_ethphy_sink_last;
wire [7:0] soc_ethphy_sink_payload_data;
wire soc_ethphy_sink_payload_last_be;
wire soc_ethphy_sink_payload_error;
wire soc_ethphy_tx_ctl_obuf;
wire [3:0] soc_ethphy_tx_data_obuf;
reg soc_ethphy_source_valid = 1'd0;
wire soc_ethphy_source_ready;
reg soc_ethphy_source_first = 1'd0;
wire soc_ethphy_source_last;
reg [7:0] soc_ethphy_source_payload_data = 8'd0;
reg soc_ethphy_source_payload_last_be = 1'd0;
reg soc_ethphy_source_payload_error = 1'd0;
wire soc_ethphy_rx_ctl_ibuf;
wire soc_ethphy_rx_ctl_idelay;
wire soc_ethphy_rx_ctl;
wire [3:0] soc_ethphy_rx_data_ibuf;
wire [3:0] soc_ethphy_rx_data_idelay;
wire [7:0] soc_ethphy_rx_data;
reg soc_ethphy_rx_ctl_d = 1'd0;
wire soc_ethphy_last;
reg [2:0] soc_ethphy_storage_full = 3'd0;
wire [2:0] soc_ethphy_storage;
reg soc_ethphy_re = 1'd0;
wire soc_ethphy_status;
wire soc_ethphy_data_w;
wire soc_ethphy_data_oe;
wire soc_ethphy_data_r;
wire soc_ethmac_tx_gap_inserter_sink_valid;
reg soc_ethmac_tx_gap_inserter_sink_ready = 1'd0;
wire soc_ethmac_tx_gap_inserter_sink_first;
wire soc_ethmac_tx_gap_inserter_sink_last;
wire [7:0] soc_ethmac_tx_gap_inserter_sink_payload_data;
wire soc_ethmac_tx_gap_inserter_sink_payload_last_be;
wire soc_ethmac_tx_gap_inserter_sink_payload_error;
reg soc_ethmac_tx_gap_inserter_source_valid = 1'd0;
wire soc_ethmac_tx_gap_inserter_source_ready;
reg soc_ethmac_tx_gap_inserter_source_first = 1'd0;
reg soc_ethmac_tx_gap_inserter_source_last = 1'd0;
reg [7:0] soc_ethmac_tx_gap_inserter_source_payload_data = 8'd0;
reg soc_ethmac_tx_gap_inserter_source_payload_last_be = 1'd0;
reg soc_ethmac_tx_gap_inserter_source_payload_error = 1'd0;
reg [3:0] soc_ethmac_tx_gap_inserter_counter = 4'd0;
reg soc_ethmac_tx_gap_inserter_counter_reset = 1'd0;
reg soc_ethmac_tx_gap_inserter_counter_ce = 1'd0;
wire soc_ethmac_rx_gap_checker_sink_valid;
reg soc_ethmac_rx_gap_checker_sink_ready = 1'd0;
wire soc_ethmac_rx_gap_checker_sink_first;
wire soc_ethmac_rx_gap_checker_sink_last;
wire [7:0] soc_ethmac_rx_gap_checker_sink_payload_data;
wire soc_ethmac_rx_gap_checker_sink_payload_last_be;
wire soc_ethmac_rx_gap_checker_sink_payload_error;
reg soc_ethmac_rx_gap_checker_source_valid = 1'd0;
wire soc_ethmac_rx_gap_checker_source_ready;
reg soc_ethmac_rx_gap_checker_source_first = 1'd0;
reg soc_ethmac_rx_gap_checker_source_last = 1'd0;
reg [7:0] soc_ethmac_rx_gap_checker_source_payload_data = 8'd0;
reg soc_ethmac_rx_gap_checker_source_payload_last_be = 1'd0;
reg soc_ethmac_rx_gap_checker_source_payload_error = 1'd0;
reg [3:0] soc_ethmac_rx_gap_checker_counter = 4'd0;
reg soc_ethmac_rx_gap_checker_counter_reset = 1'd0;
reg soc_ethmac_rx_gap_checker_counter_ce = 1'd0;
reg soc_ethmac_status = 1'd1;
wire soc_ethmac_preamble_inserter_sink_valid;
reg soc_ethmac_preamble_inserter_sink_ready = 1'd0;
wire soc_ethmac_preamble_inserter_sink_first;
wire soc_ethmac_preamble_inserter_sink_last;
wire [7:0] soc_ethmac_preamble_inserter_sink_payload_data;
wire soc_ethmac_preamble_inserter_sink_payload_last_be;
wire soc_ethmac_preamble_inserter_sink_payload_error;
reg soc_ethmac_preamble_inserter_source_valid = 1'd0;
wire soc_ethmac_preamble_inserter_source_ready;
reg soc_ethmac_preamble_inserter_source_first = 1'd0;
reg soc_ethmac_preamble_inserter_source_last = 1'd0;
reg [7:0] soc_ethmac_preamble_inserter_source_payload_data = 8'd0;
wire soc_ethmac_preamble_inserter_source_payload_last_be;
reg soc_ethmac_preamble_inserter_source_payload_error = 1'd0;
reg [63:0] soc_ethmac_preamble_inserter_preamble = 64'd15372286728091293013;
reg [2:0] soc_ethmac_preamble_inserter_cnt = 3'd0;
reg soc_ethmac_preamble_inserter_clr_cnt = 1'd0;
reg soc_ethmac_preamble_inserter_inc_cnt = 1'd0;
wire soc_ethmac_preamble_checker_sink_valid;
reg soc_ethmac_preamble_checker_sink_ready = 1'd0;
wire soc_ethmac_preamble_checker_sink_first;
wire soc_ethmac_preamble_checker_sink_last;
wire [7:0] soc_ethmac_preamble_checker_sink_payload_data;
wire soc_ethmac_preamble_checker_sink_payload_last_be;
wire soc_ethmac_preamble_checker_sink_payload_error;
reg soc_ethmac_preamble_checker_source_valid = 1'd0;
wire soc_ethmac_preamble_checker_source_ready;
reg soc_ethmac_preamble_checker_source_first = 1'd0;
reg soc_ethmac_preamble_checker_source_last = 1'd0;
wire [7:0] soc_ethmac_preamble_checker_source_payload_data;
wire soc_ethmac_preamble_checker_source_payload_last_be;
reg soc_ethmac_preamble_checker_source_payload_error = 1'd0;
reg [63:0] soc_ethmac_preamble_checker_preamble = 64'd15372286728091293013;
reg [2:0] soc_ethmac_preamble_checker_cnt = 3'd0;
reg soc_ethmac_preamble_checker_clr_cnt = 1'd0;
reg soc_ethmac_preamble_checker_inc_cnt = 1'd0;
reg soc_ethmac_preamble_checker_discard = 1'd0;
reg soc_ethmac_preamble_checker_clr_discard = 1'd0;
reg soc_ethmac_preamble_checker_set_discard = 1'd0;
reg [7:0] soc_ethmac_preamble_checker_ref = 8'd0;
wire soc_ethmac_preamble_checker_match;
wire soc_ethmac_crc32_inserter_sink_valid;
reg soc_ethmac_crc32_inserter_sink_ready = 1'd0;
wire soc_ethmac_crc32_inserter_sink_first;
wire soc_ethmac_crc32_inserter_sink_last;
wire [7:0] soc_ethmac_crc32_inserter_sink_payload_data;
wire soc_ethmac_crc32_inserter_sink_payload_last_be;
wire soc_ethmac_crc32_inserter_sink_payload_error;
reg soc_ethmac_crc32_inserter_source_valid = 1'd0;
wire soc_ethmac_crc32_inserter_source_ready;
reg soc_ethmac_crc32_inserter_source_first = 1'd0;
reg soc_ethmac_crc32_inserter_source_last = 1'd0;
reg [7:0] soc_ethmac_crc32_inserter_source_payload_data = 8'd0;
reg soc_ethmac_crc32_inserter_source_payload_last_be = 1'd0;
reg soc_ethmac_crc32_inserter_source_payload_error = 1'd0;
reg [7:0] soc_ethmac_crc32_inserter_data0 = 8'd0;
wire [31:0] soc_ethmac_crc32_inserter_value;
wire soc_ethmac_crc32_inserter_error;
wire [7:0] soc_ethmac_crc32_inserter_data1;
wire [31:0] soc_ethmac_crc32_inserter_last;
reg [31:0] soc_ethmac_crc32_inserter_next = 32'd0;
reg [31:0] soc_ethmac_crc32_inserter_reg = 32'd4294967295;
reg soc_ethmac_crc32_inserter_ce = 1'd0;
reg soc_ethmac_crc32_inserter_reset = 1'd0;
reg [1:0] soc_ethmac_crc32_inserter_cnt = 2'd3;
wire soc_ethmac_crc32_inserter_cnt_done;
reg soc_ethmac_crc32_inserter_is_ongoing0 = 1'd0;
reg soc_ethmac_crc32_inserter_is_ongoing1 = 1'd0;
wire soc_ethmac_crc32_checker_sink_sink_valid;
reg soc_ethmac_crc32_checker_sink_sink_ready = 1'd0;
wire soc_ethmac_crc32_checker_sink_sink_first;
wire soc_ethmac_crc32_checker_sink_sink_last;
wire [7:0] soc_ethmac_crc32_checker_sink_sink_payload_data;
wire soc_ethmac_crc32_checker_sink_sink_payload_last_be;
wire soc_ethmac_crc32_checker_sink_sink_payload_error;
wire soc_ethmac_crc32_checker_source_source_valid;
wire soc_ethmac_crc32_checker_source_source_ready;
reg soc_ethmac_crc32_checker_source_source_first = 1'd0;
wire soc_ethmac_crc32_checker_source_source_last;
wire [7:0] soc_ethmac_crc32_checker_source_source_payload_data;
wire soc_ethmac_crc32_checker_source_source_payload_last_be;
reg soc_ethmac_crc32_checker_source_source_payload_error = 1'd0;
wire [7:0] soc_ethmac_crc32_checker_crc_data0;
wire [31:0] soc_ethmac_crc32_checker_crc_value;
wire soc_ethmac_crc32_checker_crc_error;
wire [7:0] soc_ethmac_crc32_checker_crc_data1;
wire [31:0] soc_ethmac_crc32_checker_crc_last;
reg [31:0] soc_ethmac_crc32_checker_crc_next = 32'd0;
reg [31:0] soc_ethmac_crc32_checker_crc_reg = 32'd4294967295;
reg soc_ethmac_crc32_checker_crc_ce = 1'd0;
reg soc_ethmac_crc32_checker_crc_reset = 1'd0;
reg soc_ethmac_crc32_checker_syncfifo_sink_valid = 1'd0;
wire soc_ethmac_crc32_checker_syncfifo_sink_ready;
wire soc_ethmac_crc32_checker_syncfifo_sink_first;
wire soc_ethmac_crc32_checker_syncfifo_sink_last;
wire [7:0] soc_ethmac_crc32_checker_syncfifo_sink_payload_data;
wire soc_ethmac_crc32_checker_syncfifo_sink_payload_last_be;
wire soc_ethmac_crc32_checker_syncfifo_sink_payload_error;
wire soc_ethmac_crc32_checker_syncfifo_source_valid;
wire soc_ethmac_crc32_checker_syncfifo_source_ready;
wire soc_ethmac_crc32_checker_syncfifo_source_first;
wire soc_ethmac_crc32_checker_syncfifo_source_last;
wire [7:0] soc_ethmac_crc32_checker_syncfifo_source_payload_data;
wire soc_ethmac_crc32_checker_syncfifo_source_payload_last_be;
wire soc_ethmac_crc32_checker_syncfifo_source_payload_error;
wire soc_ethmac_crc32_checker_syncfifo_syncfifo_we;
wire soc_ethmac_crc32_checker_syncfifo_syncfifo_writable;
wire soc_ethmac_crc32_checker_syncfifo_syncfifo_re;
wire soc_ethmac_crc32_checker_syncfifo_syncfifo_readable;
wire [11:0] soc_ethmac_crc32_checker_syncfifo_syncfifo_din;
wire [11:0] soc_ethmac_crc32_checker_syncfifo_syncfifo_dout;
reg [2:0] soc_ethmac_crc32_checker_syncfifo_level = 3'd0;
reg soc_ethmac_crc32_checker_syncfifo_replace = 1'd0;
reg [2:0] soc_ethmac_crc32_checker_syncfifo_produce = 3'd0;
reg [2:0] soc_ethmac_crc32_checker_syncfifo_consume = 3'd0;
reg [2:0] soc_ethmac_crc32_checker_syncfifo_wrport_adr = 3'd0;
wire [11:0] soc_ethmac_crc32_checker_syncfifo_wrport_dat_r;
wire soc_ethmac_crc32_checker_syncfifo_wrport_we;
wire [11:0] soc_ethmac_crc32_checker_syncfifo_wrport_dat_w;
wire soc_ethmac_crc32_checker_syncfifo_do_read;
wire [2:0] soc_ethmac_crc32_checker_syncfifo_rdport_adr;
wire [11:0] soc_ethmac_crc32_checker_syncfifo_rdport_dat_r;
wire [7:0] soc_ethmac_crc32_checker_syncfifo_fifo_in_payload_data;
wire soc_ethmac_crc32_checker_syncfifo_fifo_in_payload_last_be;
wire soc_ethmac_crc32_checker_syncfifo_fifo_in_payload_error;
wire soc_ethmac_crc32_checker_syncfifo_fifo_in_first;
wire soc_ethmac_crc32_checker_syncfifo_fifo_in_last;
wire [7:0] soc_ethmac_crc32_checker_syncfifo_fifo_out_payload_data;
wire soc_ethmac_crc32_checker_syncfifo_fifo_out_payload_last_be;
wire soc_ethmac_crc32_checker_syncfifo_fifo_out_payload_error;
wire soc_ethmac_crc32_checker_syncfifo_fifo_out_first;
wire soc_ethmac_crc32_checker_syncfifo_fifo_out_last;
reg soc_ethmac_crc32_checker_fifo_reset = 1'd0;
wire soc_ethmac_crc32_checker_fifo_in;
wire soc_ethmac_crc32_checker_fifo_out;
wire soc_ethmac_crc32_checker_fifo_full;
wire soc_ethmac_padding_inserter_sink_valid;
reg soc_ethmac_padding_inserter_sink_ready = 1'd0;
wire soc_ethmac_padding_inserter_sink_first;
wire soc_ethmac_padding_inserter_sink_last;
wire [7:0] soc_ethmac_padding_inserter_sink_payload_data;
wire soc_ethmac_padding_inserter_sink_payload_last_be;
wire soc_ethmac_padding_inserter_sink_payload_error;
reg soc_ethmac_padding_inserter_source_valid = 1'd0;
wire soc_ethmac_padding_inserter_source_ready;
reg soc_ethmac_padding_inserter_source_first = 1'd0;
reg soc_ethmac_padding_inserter_source_last = 1'd0;
reg [7:0] soc_ethmac_padding_inserter_source_payload_data = 8'd0;
reg soc_ethmac_padding_inserter_source_payload_last_be = 1'd0;
reg soc_ethmac_padding_inserter_source_payload_error = 1'd0;
reg [15:0] soc_ethmac_padding_inserter_counter = 16'd1;
wire soc_ethmac_padding_inserter_counter_done;
reg soc_ethmac_padding_inserter_counter_reset = 1'd0;
reg soc_ethmac_padding_inserter_counter_ce = 1'd0;
wire soc_ethmac_padding_checker_sink_valid;
wire soc_ethmac_padding_checker_sink_ready;
wire soc_ethmac_padding_checker_sink_first;
wire soc_ethmac_padding_checker_sink_last;
wire [7:0] soc_ethmac_padding_checker_sink_payload_data;
wire soc_ethmac_padding_checker_sink_payload_last_be;
wire soc_ethmac_padding_checker_sink_payload_error;
wire soc_ethmac_padding_checker_source_valid;
wire soc_ethmac_padding_checker_source_ready;
wire soc_ethmac_padding_checker_source_first;
wire soc_ethmac_padding_checker_source_last;
wire [7:0] soc_ethmac_padding_checker_source_payload_data;
wire soc_ethmac_padding_checker_source_payload_last_be;
wire soc_ethmac_padding_checker_source_payload_error;
wire soc_ethmac_tx_last_be_sink_valid;
wire soc_ethmac_tx_last_be_sink_ready;
wire soc_ethmac_tx_last_be_sink_first;
wire soc_ethmac_tx_last_be_sink_last;
wire [7:0] soc_ethmac_tx_last_be_sink_payload_data;
wire soc_ethmac_tx_last_be_sink_payload_last_be;
wire soc_ethmac_tx_last_be_sink_payload_error;
wire soc_ethmac_tx_last_be_source_valid;
wire soc_ethmac_tx_last_be_source_ready;
reg soc_ethmac_tx_last_be_source_first = 1'd0;
wire soc_ethmac_tx_last_be_source_last;
wire [7:0] soc_ethmac_tx_last_be_source_payload_data;
reg soc_ethmac_tx_last_be_source_payload_last_be = 1'd0;
reg soc_ethmac_tx_last_be_source_payload_error = 1'd0;
reg soc_ethmac_tx_last_be_ongoing = 1'd1;
wire soc_ethmac_rx_last_be_sink_valid;
wire soc_ethmac_rx_last_be_sink_ready;
wire soc_ethmac_rx_last_be_sink_first;
wire soc_ethmac_rx_last_be_sink_last;
wire [7:0] soc_ethmac_rx_last_be_sink_payload_data;
wire soc_ethmac_rx_last_be_sink_payload_last_be;
wire soc_ethmac_rx_last_be_sink_payload_error;
wire soc_ethmac_rx_last_be_source_valid;
wire soc_ethmac_rx_last_be_source_ready;
wire soc_ethmac_rx_last_be_source_first;
wire soc_ethmac_rx_last_be_source_last;
wire [7:0] soc_ethmac_rx_last_be_source_payload_data;
reg soc_ethmac_rx_last_be_source_payload_last_be = 1'd0;
wire soc_ethmac_rx_last_be_source_payload_error;
wire soc_ethmac_tx_converter_sink_valid;
wire soc_ethmac_tx_converter_sink_ready;
wire soc_ethmac_tx_converter_sink_first;
wire soc_ethmac_tx_converter_sink_last;
wire [31:0] soc_ethmac_tx_converter_sink_payload_data;
wire [3:0] soc_ethmac_tx_converter_sink_payload_last_be;
wire [3:0] soc_ethmac_tx_converter_sink_payload_error;
wire soc_ethmac_tx_converter_source_valid;
wire soc_ethmac_tx_converter_source_ready;
wire soc_ethmac_tx_converter_source_first;
wire soc_ethmac_tx_converter_source_last;
wire [7:0] soc_ethmac_tx_converter_source_payload_data;
wire soc_ethmac_tx_converter_source_payload_last_be;
wire soc_ethmac_tx_converter_source_payload_error;
wire soc_ethmac_tx_converter_converter_sink_valid;
wire soc_ethmac_tx_converter_converter_sink_ready;
wire soc_ethmac_tx_converter_converter_sink_first;
wire soc_ethmac_tx_converter_converter_sink_last;
reg [39:0] soc_ethmac_tx_converter_converter_sink_payload_data = 40'd0;
wire soc_ethmac_tx_converter_converter_source_valid;
wire soc_ethmac_tx_converter_converter_source_ready;
wire soc_ethmac_tx_converter_converter_source_first;
wire soc_ethmac_tx_converter_converter_source_last;
reg [9:0] soc_ethmac_tx_converter_converter_source_payload_data = 10'd0;
wire soc_ethmac_tx_converter_converter_source_payload_valid_token_count;
reg [1:0] soc_ethmac_tx_converter_converter_mux = 2'd0;
wire soc_ethmac_tx_converter_converter_first;
wire soc_ethmac_tx_converter_converter_last;
wire soc_ethmac_tx_converter_source_source_valid;
wire soc_ethmac_tx_converter_source_source_ready;
wire soc_ethmac_tx_converter_source_source_first;
wire soc_ethmac_tx_converter_source_source_last;
wire [9:0] soc_ethmac_tx_converter_source_source_payload_data;
wire soc_ethmac_rx_converter_sink_valid;
wire soc_ethmac_rx_converter_sink_ready;
wire soc_ethmac_rx_converter_sink_first;
wire soc_ethmac_rx_converter_sink_last;
wire [7:0] soc_ethmac_rx_converter_sink_payload_data;
wire soc_ethmac_rx_converter_sink_payload_last_be;
wire soc_ethmac_rx_converter_sink_payload_error;
wire soc_ethmac_rx_converter_source_valid;
wire soc_ethmac_rx_converter_source_ready;
wire soc_ethmac_rx_converter_source_first;
wire soc_ethmac_rx_converter_source_last;
reg [31:0] soc_ethmac_rx_converter_source_payload_data = 32'd0;
reg [3:0] soc_ethmac_rx_converter_source_payload_last_be = 4'd0;
reg [3:0] soc_ethmac_rx_converter_source_payload_error = 4'd0;
wire soc_ethmac_rx_converter_converter_sink_valid;
wire soc_ethmac_rx_converter_converter_sink_ready;
wire soc_ethmac_rx_converter_converter_sink_first;
wire soc_ethmac_rx_converter_converter_sink_last;
wire [9:0] soc_ethmac_rx_converter_converter_sink_payload_data;
wire soc_ethmac_rx_converter_converter_source_valid;
wire soc_ethmac_rx_converter_converter_source_ready;
reg soc_ethmac_rx_converter_converter_source_first = 1'd0;
reg soc_ethmac_rx_converter_converter_source_last = 1'd0;
reg [39:0] soc_ethmac_rx_converter_converter_source_payload_data = 40'd0;
reg [2:0] soc_ethmac_rx_converter_converter_source_payload_valid_token_count = 3'd0;
reg [1:0] soc_ethmac_rx_converter_converter_demux = 2'd0;
wire soc_ethmac_rx_converter_converter_load_part;
reg soc_ethmac_rx_converter_converter_strobe_all = 1'd0;
wire soc_ethmac_rx_converter_source_source_valid;
wire soc_ethmac_rx_converter_source_source_ready;
wire soc_ethmac_rx_converter_source_source_first;
wire soc_ethmac_rx_converter_source_source_last;
wire [39:0] soc_ethmac_rx_converter_source_source_payload_data;
wire soc_ethmac_tx_cdc_sink_valid;
wire soc_ethmac_tx_cdc_sink_ready;
wire soc_ethmac_tx_cdc_sink_first;
wire soc_ethmac_tx_cdc_sink_last;
wire [31:0] soc_ethmac_tx_cdc_sink_payload_data;
wire [3:0] soc_ethmac_tx_cdc_sink_payload_last_be;
wire [3:0] soc_ethmac_tx_cdc_sink_payload_error;
wire soc_ethmac_tx_cdc_source_valid;
wire soc_ethmac_tx_cdc_source_ready;
wire soc_ethmac_tx_cdc_source_first;
wire soc_ethmac_tx_cdc_source_last;
wire [31:0] soc_ethmac_tx_cdc_source_payload_data;
wire [3:0] soc_ethmac_tx_cdc_source_payload_last_be;
wire [3:0] soc_ethmac_tx_cdc_source_payload_error;
wire soc_ethmac_tx_cdc_asyncfifo_we;
wire soc_ethmac_tx_cdc_asyncfifo_writable;
wire soc_ethmac_tx_cdc_asyncfifo_re;
wire soc_ethmac_tx_cdc_asyncfifo_readable;
wire [41:0] soc_ethmac_tx_cdc_asyncfifo_din;
wire [41:0] soc_ethmac_tx_cdc_asyncfifo_dout;
wire soc_ethmac_tx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] soc_ethmac_tx_cdc_graycounter0_q = 7'd0;
wire [6:0] soc_ethmac_tx_cdc_graycounter0_q_next;
reg [6:0] soc_ethmac_tx_cdc_graycounter0_q_binary = 7'd0;
reg [6:0] soc_ethmac_tx_cdc_graycounter0_q_next_binary = 7'd0;
wire soc_ethmac_tx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] soc_ethmac_tx_cdc_graycounter1_q = 7'd0;
wire [6:0] soc_ethmac_tx_cdc_graycounter1_q_next;
reg [6:0] soc_ethmac_tx_cdc_graycounter1_q_binary = 7'd0;
reg [6:0] soc_ethmac_tx_cdc_graycounter1_q_next_binary = 7'd0;
wire [6:0] soc_ethmac_tx_cdc_produce_rdomain;
wire [6:0] soc_ethmac_tx_cdc_consume_wdomain;
wire [5:0] soc_ethmac_tx_cdc_wrport_adr;
wire [41:0] soc_ethmac_tx_cdc_wrport_dat_r;
wire soc_ethmac_tx_cdc_wrport_we;
wire [41:0] soc_ethmac_tx_cdc_wrport_dat_w;
wire [5:0] soc_ethmac_tx_cdc_rdport_adr;
wire [41:0] soc_ethmac_tx_cdc_rdport_dat_r;
wire [31:0] soc_ethmac_tx_cdc_fifo_in_payload_data;
wire [3:0] soc_ethmac_tx_cdc_fifo_in_payload_last_be;
wire [3:0] soc_ethmac_tx_cdc_fifo_in_payload_error;
wire soc_ethmac_tx_cdc_fifo_in_first;
wire soc_ethmac_tx_cdc_fifo_in_last;
wire [31:0] soc_ethmac_tx_cdc_fifo_out_payload_data;
wire [3:0] soc_ethmac_tx_cdc_fifo_out_payload_last_be;
wire [3:0] soc_ethmac_tx_cdc_fifo_out_payload_error;
wire soc_ethmac_tx_cdc_fifo_out_first;
wire soc_ethmac_tx_cdc_fifo_out_last;
wire soc_ethmac_rx_cdc_sink_valid;
wire soc_ethmac_rx_cdc_sink_ready;
wire soc_ethmac_rx_cdc_sink_first;
wire soc_ethmac_rx_cdc_sink_last;
wire [31:0] soc_ethmac_rx_cdc_sink_payload_data;
wire [3:0] soc_ethmac_rx_cdc_sink_payload_last_be;
wire [3:0] soc_ethmac_rx_cdc_sink_payload_error;
wire soc_ethmac_rx_cdc_source_valid;
wire soc_ethmac_rx_cdc_source_ready;
wire soc_ethmac_rx_cdc_source_first;
wire soc_ethmac_rx_cdc_source_last;
wire [31:0] soc_ethmac_rx_cdc_source_payload_data;
wire [3:0] soc_ethmac_rx_cdc_source_payload_last_be;
wire [3:0] soc_ethmac_rx_cdc_source_payload_error;
wire soc_ethmac_rx_cdc_asyncfifo_we;
wire soc_ethmac_rx_cdc_asyncfifo_writable;
wire soc_ethmac_rx_cdc_asyncfifo_re;
wire soc_ethmac_rx_cdc_asyncfifo_readable;
wire [41:0] soc_ethmac_rx_cdc_asyncfifo_din;
wire [41:0] soc_ethmac_rx_cdc_asyncfifo_dout;
wire soc_ethmac_rx_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [6:0] soc_ethmac_rx_cdc_graycounter0_q = 7'd0;
wire [6:0] soc_ethmac_rx_cdc_graycounter0_q_next;
reg [6:0] soc_ethmac_rx_cdc_graycounter0_q_binary = 7'd0;
reg [6:0] soc_ethmac_rx_cdc_graycounter0_q_next_binary = 7'd0;
wire soc_ethmac_rx_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [6:0] soc_ethmac_rx_cdc_graycounter1_q = 7'd0;
wire [6:0] soc_ethmac_rx_cdc_graycounter1_q_next;
reg [6:0] soc_ethmac_rx_cdc_graycounter1_q_binary = 7'd0;
reg [6:0] soc_ethmac_rx_cdc_graycounter1_q_next_binary = 7'd0;
wire [6:0] soc_ethmac_rx_cdc_produce_rdomain;
wire [6:0] soc_ethmac_rx_cdc_consume_wdomain;
wire [5:0] soc_ethmac_rx_cdc_wrport_adr;
wire [41:0] soc_ethmac_rx_cdc_wrport_dat_r;
wire soc_ethmac_rx_cdc_wrport_we;
wire [41:0] soc_ethmac_rx_cdc_wrport_dat_w;
wire [5:0] soc_ethmac_rx_cdc_rdport_adr;
wire [41:0] soc_ethmac_rx_cdc_rdport_dat_r;
wire [31:0] soc_ethmac_rx_cdc_fifo_in_payload_data;
wire [3:0] soc_ethmac_rx_cdc_fifo_in_payload_last_be;
wire [3:0] soc_ethmac_rx_cdc_fifo_in_payload_error;
wire soc_ethmac_rx_cdc_fifo_in_first;
wire soc_ethmac_rx_cdc_fifo_in_last;
wire [31:0] soc_ethmac_rx_cdc_fifo_out_payload_data;
wire [3:0] soc_ethmac_rx_cdc_fifo_out_payload_last_be;
wire [3:0] soc_ethmac_rx_cdc_fifo_out_payload_error;
wire soc_ethmac_rx_cdc_fifo_out_first;
wire soc_ethmac_rx_cdc_fifo_out_last;
wire soc_ethmac_sink_valid;
wire soc_ethmac_sink_ready;
wire soc_ethmac_sink_first;
wire soc_ethmac_sink_last;
wire [31:0] soc_ethmac_sink_payload_data;
wire [3:0] soc_ethmac_sink_payload_last_be;
wire [3:0] soc_ethmac_sink_payload_error;
wire soc_ethmac_source_valid;
wire soc_ethmac_source_ready;
wire soc_ethmac_source_first;
wire soc_ethmac_source_last;
wire [31:0] soc_ethmac_source_payload_data;
wire [3:0] soc_ethmac_source_payload_last_be;
wire [3:0] soc_ethmac_source_payload_error;
wire [29:0] soc_ethmac_bus_adr;
wire [31:0] soc_ethmac_bus_dat_w;
wire [31:0] soc_ethmac_bus_dat_r;
wire [3:0] soc_ethmac_bus_sel;
wire soc_ethmac_bus_cyc;
wire soc_ethmac_bus_stb;
wire soc_ethmac_bus_ack;
wire soc_ethmac_bus_we;
wire [2:0] soc_ethmac_bus_cti;
wire [1:0] soc_ethmac_bus_bte;
wire soc_ethmac_bus_err;
wire soc_ethmac_writer_sink_sink_valid;
reg soc_ethmac_writer_sink_sink_ready = 1'd1;
wire soc_ethmac_writer_sink_sink_first;
wire soc_ethmac_writer_sink_sink_last;
wire [31:0] soc_ethmac_writer_sink_sink_payload_data;
wire [3:0] soc_ethmac_writer_sink_sink_payload_last_be;
wire [3:0] soc_ethmac_writer_sink_sink_payload_error;
wire soc_ethmac_writer_slot_status;
wire [31:0] soc_ethmac_writer_length_status;
wire soc_ethmac_writer_irq;
wire soc_ethmac_writer_available_status;
wire soc_ethmac_writer_available_pending;
wire soc_ethmac_writer_available_trigger;
reg soc_ethmac_writer_available_clear = 1'd0;
wire soc_ethmac_writer_status_re;
wire soc_ethmac_writer_status_r;
wire soc_ethmac_writer_status_w;
wire soc_ethmac_writer_pending_re;
wire soc_ethmac_writer_pending_r;
wire soc_ethmac_writer_pending_w;
reg soc_ethmac_writer_storage_full = 1'd0;
wire soc_ethmac_writer_storage;
reg soc_ethmac_writer_re = 1'd0;
reg [2:0] soc_ethmac_writer_increment = 3'd0;
reg [31:0] soc_ethmac_writer_counter = 32'd0;
reg soc_ethmac_writer_counter_reset = 1'd0;
reg soc_ethmac_writer_counter_ce = 1'd0;
reg soc_ethmac_writer_slot = 1'd0;
reg soc_ethmac_writer_slot_ce = 1'd0;
reg soc_ethmac_writer_ongoing = 1'd0;
reg soc_ethmac_writer_fifo_sink_valid = 1'd0;
wire soc_ethmac_writer_fifo_sink_ready;
reg soc_ethmac_writer_fifo_sink_first = 1'd0;
reg soc_ethmac_writer_fifo_sink_last = 1'd0;
wire soc_ethmac_writer_fifo_sink_payload_slot;
wire [31:0] soc_ethmac_writer_fifo_sink_payload_length;
wire soc_ethmac_writer_fifo_source_valid;
wire soc_ethmac_writer_fifo_source_ready;
wire soc_ethmac_writer_fifo_source_first;
wire soc_ethmac_writer_fifo_source_last;
wire soc_ethmac_writer_fifo_source_payload_slot;
wire [31:0] soc_ethmac_writer_fifo_source_payload_length;
wire soc_ethmac_writer_fifo_syncfifo_we;
wire soc_ethmac_writer_fifo_syncfifo_writable;
wire soc_ethmac_writer_fifo_syncfifo_re;
wire soc_ethmac_writer_fifo_syncfifo_readable;
wire [34:0] soc_ethmac_writer_fifo_syncfifo_din;
wire [34:0] soc_ethmac_writer_fifo_syncfifo_dout;
reg [1:0] soc_ethmac_writer_fifo_level = 2'd0;
reg soc_ethmac_writer_fifo_replace = 1'd0;
reg soc_ethmac_writer_fifo_produce = 1'd0;
reg soc_ethmac_writer_fifo_consume = 1'd0;
reg soc_ethmac_writer_fifo_wrport_adr = 1'd0;
wire [34:0] soc_ethmac_writer_fifo_wrport_dat_r;
wire soc_ethmac_writer_fifo_wrport_we;
wire [34:0] soc_ethmac_writer_fifo_wrport_dat_w;
wire soc_ethmac_writer_fifo_do_read;
wire soc_ethmac_writer_fifo_rdport_adr;
wire [34:0] soc_ethmac_writer_fifo_rdport_dat_r;
wire soc_ethmac_writer_fifo_fifo_in_payload_slot;
wire [31:0] soc_ethmac_writer_fifo_fifo_in_payload_length;
wire soc_ethmac_writer_fifo_fifo_in_first;
wire soc_ethmac_writer_fifo_fifo_in_last;
wire soc_ethmac_writer_fifo_fifo_out_payload_slot;
wire [31:0] soc_ethmac_writer_fifo_fifo_out_payload_length;
wire soc_ethmac_writer_fifo_fifo_out_first;
wire soc_ethmac_writer_fifo_fifo_out_last;
reg [8:0] soc_ethmac_writer_memory0_adr = 9'd0;
wire [31:0] soc_ethmac_writer_memory0_dat_r;
reg soc_ethmac_writer_memory0_we = 1'd0;
reg [31:0] soc_ethmac_writer_memory0_dat_w = 32'd0;
reg [8:0] soc_ethmac_writer_memory1_adr = 9'd0;
wire [31:0] soc_ethmac_writer_memory1_dat_r;
reg soc_ethmac_writer_memory1_we = 1'd0;
reg [31:0] soc_ethmac_writer_memory1_dat_w = 32'd0;
reg soc_ethmac_reader_source_source_valid = 1'd0;
wire soc_ethmac_reader_source_source_ready;
reg soc_ethmac_reader_source_source_first = 1'd0;
reg soc_ethmac_reader_source_source_last = 1'd0;
reg [31:0] soc_ethmac_reader_source_source_payload_data = 32'd0;
reg [3:0] soc_ethmac_reader_source_source_payload_last_be = 4'd0;
reg [3:0] soc_ethmac_reader_source_source_payload_error = 4'd0;
wire soc_ethmac_reader_start_re;
wire soc_ethmac_reader_start_r;
reg soc_ethmac_reader_start_w = 1'd0;
wire soc_ethmac_reader_ready_status;
reg soc_ethmac_reader_slot_storage_full = 1'd0;
wire soc_ethmac_reader_slot_storage;
reg soc_ethmac_reader_slot_re = 1'd0;
reg [10:0] soc_ethmac_reader_length_storage_full = 11'd0;
wire [10:0] soc_ethmac_reader_length_storage;
reg soc_ethmac_reader_length_re = 1'd0;
wire soc_ethmac_reader_irq;
wire soc_ethmac_reader_done_status;
reg soc_ethmac_reader_done_pending = 1'd0;
reg soc_ethmac_reader_done_trigger = 1'd0;
reg soc_ethmac_reader_done_clear = 1'd0;
wire soc_ethmac_reader_eventmanager_status_re;
wire soc_ethmac_reader_eventmanager_status_r;
wire soc_ethmac_reader_eventmanager_status_w;
wire soc_ethmac_reader_eventmanager_pending_re;
wire soc_ethmac_reader_eventmanager_pending_r;
wire soc_ethmac_reader_eventmanager_pending_w;
reg soc_ethmac_reader_eventmanager_storage_full = 1'd0;
wire soc_ethmac_reader_eventmanager_storage;
reg soc_ethmac_reader_eventmanager_re = 1'd0;
wire soc_ethmac_reader_fifo_sink_valid;
wire soc_ethmac_reader_fifo_sink_ready;
reg soc_ethmac_reader_fifo_sink_first = 1'd0;
reg soc_ethmac_reader_fifo_sink_last = 1'd0;
wire soc_ethmac_reader_fifo_sink_payload_slot;
wire [10:0] soc_ethmac_reader_fifo_sink_payload_length;
wire soc_ethmac_reader_fifo_source_valid;
reg soc_ethmac_reader_fifo_source_ready = 1'd0;
wire soc_ethmac_reader_fifo_source_first;
wire soc_ethmac_reader_fifo_source_last;
wire soc_ethmac_reader_fifo_source_payload_slot;
wire [10:0] soc_ethmac_reader_fifo_source_payload_length;
wire soc_ethmac_reader_fifo_syncfifo_we;
wire soc_ethmac_reader_fifo_syncfifo_writable;
wire soc_ethmac_reader_fifo_syncfifo_re;
wire soc_ethmac_reader_fifo_syncfifo_readable;
wire [13:0] soc_ethmac_reader_fifo_syncfifo_din;
wire [13:0] soc_ethmac_reader_fifo_syncfifo_dout;
reg [1:0] soc_ethmac_reader_fifo_level = 2'd0;
reg soc_ethmac_reader_fifo_replace = 1'd0;
reg soc_ethmac_reader_fifo_produce = 1'd0;
reg soc_ethmac_reader_fifo_consume = 1'd0;
reg soc_ethmac_reader_fifo_wrport_adr = 1'd0;
wire [13:0] soc_ethmac_reader_fifo_wrport_dat_r;
wire soc_ethmac_reader_fifo_wrport_we;
wire [13:0] soc_ethmac_reader_fifo_wrport_dat_w;
wire soc_ethmac_reader_fifo_do_read;
wire soc_ethmac_reader_fifo_rdport_adr;
wire [13:0] soc_ethmac_reader_fifo_rdport_dat_r;
wire soc_ethmac_reader_fifo_fifo_in_payload_slot;
wire [10:0] soc_ethmac_reader_fifo_fifo_in_payload_length;
wire soc_ethmac_reader_fifo_fifo_in_first;
wire soc_ethmac_reader_fifo_fifo_in_last;
wire soc_ethmac_reader_fifo_fifo_out_payload_slot;
wire [10:0] soc_ethmac_reader_fifo_fifo_out_payload_length;
wire soc_ethmac_reader_fifo_fifo_out_first;
wire soc_ethmac_reader_fifo_fifo_out_last;
reg [10:0] soc_ethmac_reader_counter = 11'd0;
reg soc_ethmac_reader_counter_reset = 1'd0;
reg soc_ethmac_reader_counter_ce = 1'd0;
wire soc_ethmac_reader_last;
wire [8:0] soc_ethmac_reader_memory0_adr;
wire [31:0] soc_ethmac_reader_memory0_dat_r;
wire [8:0] soc_ethmac_reader_memory1_adr;
wire [31:0] soc_ethmac_reader_memory1_dat_r;
wire soc_ethmac_ev_irq;
wire [29:0] soc_ethmac_sram0_bus_adr0;
wire [31:0] soc_ethmac_sram0_bus_dat_w0;
wire [31:0] soc_ethmac_sram0_bus_dat_r0;
wire [3:0] soc_ethmac_sram0_bus_sel0;
wire soc_ethmac_sram0_bus_cyc0;
wire soc_ethmac_sram0_bus_stb0;
reg soc_ethmac_sram0_bus_ack0 = 1'd0;
wire soc_ethmac_sram0_bus_we0;
wire [2:0] soc_ethmac_sram0_bus_cti0;
wire [1:0] soc_ethmac_sram0_bus_bte0;
reg soc_ethmac_sram0_bus_err0 = 1'd0;
wire [8:0] soc_ethmac_sram0_adr0;
wire [31:0] soc_ethmac_sram0_dat_r0;
wire [29:0] soc_ethmac_sram1_bus_adr0;
wire [31:0] soc_ethmac_sram1_bus_dat_w0;
wire [31:0] soc_ethmac_sram1_bus_dat_r0;
wire [3:0] soc_ethmac_sram1_bus_sel0;
wire soc_ethmac_sram1_bus_cyc0;
wire soc_ethmac_sram1_bus_stb0;
reg soc_ethmac_sram1_bus_ack0 = 1'd0;
wire soc_ethmac_sram1_bus_we0;
wire [2:0] soc_ethmac_sram1_bus_cti0;
wire [1:0] soc_ethmac_sram1_bus_bte0;
reg soc_ethmac_sram1_bus_err0 = 1'd0;
wire [8:0] soc_ethmac_sram1_adr0;
wire [31:0] soc_ethmac_sram1_dat_r0;
wire [29:0] soc_ethmac_sram0_bus_adr1;
wire [31:0] soc_ethmac_sram0_bus_dat_w1;
wire [31:0] soc_ethmac_sram0_bus_dat_r1;
wire [3:0] soc_ethmac_sram0_bus_sel1;
wire soc_ethmac_sram0_bus_cyc1;
wire soc_ethmac_sram0_bus_stb1;
reg soc_ethmac_sram0_bus_ack1 = 1'd0;
wire soc_ethmac_sram0_bus_we1;
wire [2:0] soc_ethmac_sram0_bus_cti1;
wire [1:0] soc_ethmac_sram0_bus_bte1;
reg soc_ethmac_sram0_bus_err1 = 1'd0;
wire [8:0] soc_ethmac_sram0_adr1;
wire [31:0] soc_ethmac_sram0_dat_r1;
reg [3:0] soc_ethmac_sram0_we = 4'd0;
wire [31:0] soc_ethmac_sram0_dat_w;
wire [29:0] soc_ethmac_sram1_bus_adr1;
wire [31:0] soc_ethmac_sram1_bus_dat_w1;
wire [31:0] soc_ethmac_sram1_bus_dat_r1;
wire [3:0] soc_ethmac_sram1_bus_sel1;
wire soc_ethmac_sram1_bus_cyc1;
wire soc_ethmac_sram1_bus_stb1;
reg soc_ethmac_sram1_bus_ack1 = 1'd0;
wire soc_ethmac_sram1_bus_we1;
wire [2:0] soc_ethmac_sram1_bus_cti1;
wire [1:0] soc_ethmac_sram1_bus_bte1;
reg soc_ethmac_sram1_bus_err1 = 1'd0;
wire [8:0] soc_ethmac_sram1_adr1;
wire [31:0] soc_ethmac_sram1_dat_r1;
reg [3:0] soc_ethmac_sram1_we = 4'd0;
wire [31:0] soc_ethmac_sram1_dat_w;
reg [3:0] soc_ethmac_slave_sel = 4'd0;
reg [3:0] soc_ethmac_slave_sel_r = 4'd0;
wire soc_litedramcrossbar_cmd_valid;
wire soc_litedramcrossbar_cmd_ready;
wire soc_litedramcrossbar_cmd_payload_we;
wire [24:0] soc_litedramcrossbar_cmd_payload_adr;
wire soc_litedramcrossbar_wdata_valid;
wire soc_litedramcrossbar_wdata_ready;
wire [127:0] soc_litedramcrossbar_wdata_payload_data;
wire [15:0] soc_litedramcrossbar_wdata_payload_we;
wire soc_litedramcrossbar_rdata_valid;
wire [127:0] soc_litedramcrossbar_rdata_payload_data;
wire soc_edid_status;
reg soc_edid_storage_full = 1'd0;
wire soc_edid_storage;
reg soc_edid_re = 1'd0;
wire soc_edid_scl_raw;
reg soc_edid_sda_i = 1'd0;
wire soc_edid_sda_raw;
reg soc_edid_sda_drv = 1'd0;
reg soc_edid_sda_drv_reg = 1'd0;
wire soc_edid_sda_i_async;
wire soc_edid_sda_o;
reg soc_edid_scl_i = 1'd0;
reg [5:0] soc_edid_samp_count = 6'd0;
reg soc_edid_samp_carry = 1'd0;
reg soc_edid_scl_r = 1'd0;
reg soc_edid_sda_r = 1'd0;
wire soc_edid_scl_rising;
wire soc_edid_sda_rising;
wire soc_edid_sda_falling;
wire soc_edid_start;
reg [7:0] soc_edid_din = 8'd0;
reg [3:0] soc_edid_counter = 4'd0;
reg soc_edid_is_read = 1'd0;
reg soc_edid_update_is_read = 1'd0;
reg [6:0] soc_edid_offset_counter = 7'd0;
reg soc_edid_oc_load = 1'd0;
reg soc_edid_oc_inc = 1'd0;
wire [6:0] soc_edid_adr;
wire [7:0] soc_edid_dat_r;
reg soc_edid_data_bit = 1'd0;
reg soc_edid_zero_drv = 1'd0;
reg soc_edid_data_drv = 1'd0;
reg soc_edid_data_drv_en = 1'd0;
reg soc_edid_data_drv_stop = 1'd0;
reg soc_mmcm_reset_storage_full = 1'd1;
wire soc_mmcm_reset_storage;
reg soc_mmcm_reset_re = 1'd0;
wire soc_locked_status;
wire soc_mmcm_read_re;
wire soc_mmcm_read_r;
reg soc_mmcm_read_w = 1'd0;
wire soc_mmcm_write_re;
wire soc_mmcm_write_r;
reg soc_mmcm_write_w = 1'd0;
reg soc_mmcm_drdy_status = 1'd0;
reg [6:0] soc_mmcm_adr_storage_full = 7'd0;
wire [6:0] soc_mmcm_adr_storage;
reg soc_mmcm_adr_re = 1'd0;
reg [15:0] soc_mmcm_dat_w_storage_full = 16'd0;
wire [15:0] soc_mmcm_dat_w_storage;
reg soc_mmcm_dat_w_re = 1'd0;
wire [15:0] soc_mmcm_dat_r_status;
wire soc_locked;
wire hdmi_in0_pix_clk;
wire hdmi_in0_pix_rst;
wire pix1p25x_clk;
wire pix1p25x_rst;
wire hdmi_in0_pix5x_clk;
wire soc_clk_input;
wire soc_clk_input_bufg;
wire soc_mmcm_fb;
wire soc_mmcm_locked;
wire soc_mmcm_clk0;
wire soc_mmcm_clk1;
wire soc_mmcm_clk2;
wire soc_mmcm_drdy;
wire [9:0] soc_s7datacapture0_d;
wire soc_s7datacapture0_dly_ctl_re;
wire [4:0] soc_s7datacapture0_dly_ctl_r;
reg [4:0] soc_s7datacapture0_dly_ctl_w = 5'd0;
wire [1:0] soc_s7datacapture0_status;
wire soc_s7datacapture0_phase_reset_re;
wire soc_s7datacapture0_phase_reset_r;
reg soc_s7datacapture0_phase_reset_w = 1'd0;
wire soc_s7datacapture0_serdes_m_i_nodelay;
wire soc_s7datacapture0_serdes_s_i_nodelay;
wire soc_s7datacapture0_delay_rst;
wire soc_s7datacapture0_delay_master_inc;
wire soc_s7datacapture0_delay_master_ce;
wire soc_s7datacapture0_delay_slave_inc;
wire soc_s7datacapture0_delay_slave_ce;
wire soc_s7datacapture0_serdes_m_i_delayed;
wire [7:0] soc_s7datacapture0_serdes_m_q;
wire [7:0] soc_s7datacapture0_serdes_m_d;
wire soc_s7datacapture0_serdes_s_i_delayed;
wire [7:0] soc_s7datacapture0_serdes_s_q;
wire [7:0] soc_s7datacapture0_serdes_s_d;
wire [7:0] soc_s7datacapture0_gearbox_i;
reg [9:0] soc_s7datacapture0_gearbox_o = 10'd0;
wire soc_s7datacapture0_gearbox_rst;
wire data0_cap_write_clk;
wire data0_cap_write_rst;
wire data0_cap_read_clk;
wire data0_cap_read_rst;
reg [79:0] soc_s7datacapture0_gearbox_storage = 80'd0;
reg [3:0] soc_s7datacapture0_gearbox_wrpointer = 4'd5;
reg [2:0] soc_s7datacapture0_gearbox_rdpointer = 3'd0;
wire [7:0] soc_s7datacapture0_mdata;
wire [7:0] soc_s7datacapture0_sdata;
wire soc_s7datacapture0_inc;
wire soc_s7datacapture0_dec;
wire soc_s7datacapture0_transition;
reg [7:0] soc_s7datacapture0_mdata_d = 8'd0;
reg [7:0] soc_s7datacapture0_lateness = 8'd128;
wire soc_s7datacapture0_too_late;
wire soc_s7datacapture0_too_early;
wire soc_s7datacapture0_reset_lateness;
wire soc_s7datacapture0_do_delay_rst_i;
wire soc_s7datacapture0_do_delay_rst_o;
reg soc_s7datacapture0_do_delay_rst_toggle_i = 1'd0;
wire soc_s7datacapture0_do_delay_rst_toggle_o;
reg soc_s7datacapture0_do_delay_rst_toggle_o_r = 1'd0;
wire soc_s7datacapture0_do_delay_master_inc_i;
wire soc_s7datacapture0_do_delay_master_inc_o;
reg soc_s7datacapture0_do_delay_master_inc_toggle_i = 1'd0;
wire soc_s7datacapture0_do_delay_master_inc_toggle_o;
reg soc_s7datacapture0_do_delay_master_inc_toggle_o_r = 1'd0;
wire soc_s7datacapture0_do_delay_master_dec_i;
wire soc_s7datacapture0_do_delay_master_dec_o;
reg soc_s7datacapture0_do_delay_master_dec_toggle_i = 1'd0;
wire soc_s7datacapture0_do_delay_master_dec_toggle_o;
reg soc_s7datacapture0_do_delay_master_dec_toggle_o_r = 1'd0;
wire soc_s7datacapture0_do_delay_slave_inc_i;
wire soc_s7datacapture0_do_delay_slave_inc_o;
reg soc_s7datacapture0_do_delay_slave_inc_toggle_i = 1'd0;
wire soc_s7datacapture0_do_delay_slave_inc_toggle_o;
reg soc_s7datacapture0_do_delay_slave_inc_toggle_o_r = 1'd0;
wire soc_s7datacapture0_do_delay_slave_dec_i;
wire soc_s7datacapture0_do_delay_slave_dec_o;
reg soc_s7datacapture0_do_delay_slave_dec_toggle_i = 1'd0;
wire soc_s7datacapture0_do_delay_slave_dec_toggle_o;
reg soc_s7datacapture0_do_delay_slave_dec_toggle_o_r = 1'd0;
wire soc_s7datacapture0_do_reset_lateness_i;
wire soc_s7datacapture0_do_reset_lateness_o;
reg soc_s7datacapture0_do_reset_lateness_toggle_i = 1'd0;
wire soc_s7datacapture0_do_reset_lateness_toggle_o;
reg soc_s7datacapture0_do_reset_lateness_toggle_o_r = 1'd0;
wire [9:0] soc_charsync0_raw_data;
reg soc_charsync0_synced = 1'd0;
reg [9:0] soc_charsync0_data = 10'd0;
wire soc_charsync0_char_synced_status;
wire [3:0] soc_charsync0_ctl_pos_status;
reg [9:0] soc_charsync0_raw_data1 = 10'd0;
wire [19:0] soc_charsync0_raw;
reg soc_charsync0_found_control = 1'd0;
reg [3:0] soc_charsync0_control_position = 4'd0;
reg [2:0] soc_charsync0_control_counter = 3'd0;
reg [3:0] soc_charsync0_previous_control_position = 4'd0;
reg [3:0] soc_charsync0_word_sel = 4'd0;
wire [9:0] soc_wer0_data;
wire soc_wer0_update_re;
wire soc_wer0_update_r;
reg soc_wer0_update_w = 1'd0;
reg [23:0] soc_wer0_status = 24'd0;
reg [8:0] soc_wer0_data_r = 9'd0;
reg [7:0] soc_wer0_transitions = 8'd0;
reg [3:0] soc_wer0_transition_count = 4'd0;
reg soc_wer0_is_control = 1'd0;
reg soc_wer0_is_error = 1'd0;
reg [23:0] soc_wer0_period_counter = 24'd0;
reg soc_wer0_period_done = 1'd0;
reg [23:0] soc_wer0_wer_counter = 24'd0;
reg [23:0] soc_wer0_wer_counter_r = 24'd0;
reg soc_wer0_wer_counter_r_updated = 1'd0;
reg [23:0] soc_wer0_wer_counter_sys = 24'd0;
wire soc_wer0_i;
wire soc_wer0_o;
reg soc_wer0_toggle_i = 1'd0;
wire soc_wer0_toggle_o;
reg soc_wer0_toggle_o_r = 1'd0;
wire soc_decoding0_valid_i;
wire [9:0] soc_decoding0_input;
reg soc_decoding0_valid_o = 1'd0;
reg [7:0] soc_decoding0_output_d = 8'd0;
reg [1:0] soc_decoding0_output_c = 2'd0;
reg soc_decoding0_output_de = 1'd0;
wire [9:0] soc_s7datacapture1_d;
wire soc_s7datacapture1_dly_ctl_re;
wire [4:0] soc_s7datacapture1_dly_ctl_r;
reg [4:0] soc_s7datacapture1_dly_ctl_w = 5'd0;
wire [1:0] soc_s7datacapture1_status;
wire soc_s7datacapture1_phase_reset_re;
wire soc_s7datacapture1_phase_reset_r;
reg soc_s7datacapture1_phase_reset_w = 1'd0;
wire soc_s7datacapture1_serdes_m_i_nodelay;
wire soc_s7datacapture1_serdes_s_i_nodelay;
wire soc_s7datacapture1_delay_rst;
wire soc_s7datacapture1_delay_master_inc;
wire soc_s7datacapture1_delay_master_ce;
wire soc_s7datacapture1_delay_slave_inc;
wire soc_s7datacapture1_delay_slave_ce;
wire soc_s7datacapture1_serdes_m_i_delayed;
wire [7:0] soc_s7datacapture1_serdes_m_q;
wire [7:0] soc_s7datacapture1_serdes_m_d;
wire soc_s7datacapture1_serdes_s_i_delayed;
wire [7:0] soc_s7datacapture1_serdes_s_q;
wire [7:0] soc_s7datacapture1_serdes_s_d;
wire [7:0] soc_s7datacapture1_gearbox_i;
reg [9:0] soc_s7datacapture1_gearbox_o = 10'd0;
wire soc_s7datacapture1_gearbox_rst;
wire data1_cap_write_clk;
wire data1_cap_write_rst;
wire data1_cap_read_clk;
wire data1_cap_read_rst;
reg [79:0] soc_s7datacapture1_gearbox_storage = 80'd0;
reg [3:0] soc_s7datacapture1_gearbox_wrpointer = 4'd5;
reg [2:0] soc_s7datacapture1_gearbox_rdpointer = 3'd0;
wire [7:0] soc_s7datacapture1_mdata;
wire [7:0] soc_s7datacapture1_sdata;
wire soc_s7datacapture1_inc;
wire soc_s7datacapture1_dec;
wire soc_s7datacapture1_transition;
reg [7:0] soc_s7datacapture1_mdata_d = 8'd0;
reg [7:0] soc_s7datacapture1_lateness = 8'd128;
wire soc_s7datacapture1_too_late;
wire soc_s7datacapture1_too_early;
wire soc_s7datacapture1_reset_lateness;
wire soc_s7datacapture1_do_delay_rst_i;
wire soc_s7datacapture1_do_delay_rst_o;
reg soc_s7datacapture1_do_delay_rst_toggle_i = 1'd0;
wire soc_s7datacapture1_do_delay_rst_toggle_o;
reg soc_s7datacapture1_do_delay_rst_toggle_o_r = 1'd0;
wire soc_s7datacapture1_do_delay_master_inc_i;
wire soc_s7datacapture1_do_delay_master_inc_o;
reg soc_s7datacapture1_do_delay_master_inc_toggle_i = 1'd0;
wire soc_s7datacapture1_do_delay_master_inc_toggle_o;
reg soc_s7datacapture1_do_delay_master_inc_toggle_o_r = 1'd0;
wire soc_s7datacapture1_do_delay_master_dec_i;
wire soc_s7datacapture1_do_delay_master_dec_o;
reg soc_s7datacapture1_do_delay_master_dec_toggle_i = 1'd0;
wire soc_s7datacapture1_do_delay_master_dec_toggle_o;
reg soc_s7datacapture1_do_delay_master_dec_toggle_o_r = 1'd0;
wire soc_s7datacapture1_do_delay_slave_inc_i;
wire soc_s7datacapture1_do_delay_slave_inc_o;
reg soc_s7datacapture1_do_delay_slave_inc_toggle_i = 1'd0;
wire soc_s7datacapture1_do_delay_slave_inc_toggle_o;
reg soc_s7datacapture1_do_delay_slave_inc_toggle_o_r = 1'd0;
wire soc_s7datacapture1_do_delay_slave_dec_i;
wire soc_s7datacapture1_do_delay_slave_dec_o;
reg soc_s7datacapture1_do_delay_slave_dec_toggle_i = 1'd0;
wire soc_s7datacapture1_do_delay_slave_dec_toggle_o;
reg soc_s7datacapture1_do_delay_slave_dec_toggle_o_r = 1'd0;
wire soc_s7datacapture1_do_reset_lateness_i;
wire soc_s7datacapture1_do_reset_lateness_o;
reg soc_s7datacapture1_do_reset_lateness_toggle_i = 1'd0;
wire soc_s7datacapture1_do_reset_lateness_toggle_o;
reg soc_s7datacapture1_do_reset_lateness_toggle_o_r = 1'd0;
wire [9:0] soc_charsync1_raw_data;
reg soc_charsync1_synced = 1'd0;
reg [9:0] soc_charsync1_data = 10'd0;
wire soc_charsync1_char_synced_status;
wire [3:0] soc_charsync1_ctl_pos_status;
reg [9:0] soc_charsync1_raw_data1 = 10'd0;
wire [19:0] soc_charsync1_raw;
reg soc_charsync1_found_control = 1'd0;
reg [3:0] soc_charsync1_control_position = 4'd0;
reg [2:0] soc_charsync1_control_counter = 3'd0;
reg [3:0] soc_charsync1_previous_control_position = 4'd0;
reg [3:0] soc_charsync1_word_sel = 4'd0;
wire [9:0] soc_wer1_data;
wire soc_wer1_update_re;
wire soc_wer1_update_r;
reg soc_wer1_update_w = 1'd0;
reg [23:0] soc_wer1_status = 24'd0;
reg [8:0] soc_wer1_data_r = 9'd0;
reg [7:0] soc_wer1_transitions = 8'd0;
reg [3:0] soc_wer1_transition_count = 4'd0;
reg soc_wer1_is_control = 1'd0;
reg soc_wer1_is_error = 1'd0;
reg [23:0] soc_wer1_period_counter = 24'd0;
reg soc_wer1_period_done = 1'd0;
reg [23:0] soc_wer1_wer_counter = 24'd0;
reg [23:0] soc_wer1_wer_counter_r = 24'd0;
reg soc_wer1_wer_counter_r_updated = 1'd0;
reg [23:0] soc_wer1_wer_counter_sys = 24'd0;
wire soc_wer1_i;
wire soc_wer1_o;
reg soc_wer1_toggle_i = 1'd0;
wire soc_wer1_toggle_o;
reg soc_wer1_toggle_o_r = 1'd0;
wire soc_decoding1_valid_i;
wire [9:0] soc_decoding1_input;
reg soc_decoding1_valid_o = 1'd0;
reg [7:0] soc_decoding1_output_d = 8'd0;
reg [1:0] soc_decoding1_output_c = 2'd0;
reg soc_decoding1_output_de = 1'd0;
wire [9:0] soc_s7datacapture2_d;
wire soc_s7datacapture2_dly_ctl_re;
wire [4:0] soc_s7datacapture2_dly_ctl_r;
reg [4:0] soc_s7datacapture2_dly_ctl_w = 5'd0;
wire [1:0] soc_s7datacapture2_status;
wire soc_s7datacapture2_phase_reset_re;
wire soc_s7datacapture2_phase_reset_r;
reg soc_s7datacapture2_phase_reset_w = 1'd0;
wire soc_s7datacapture2_serdes_m_i_nodelay;
wire soc_s7datacapture2_serdes_s_i_nodelay;
wire soc_s7datacapture2_delay_rst;
wire soc_s7datacapture2_delay_master_inc;
wire soc_s7datacapture2_delay_master_ce;
wire soc_s7datacapture2_delay_slave_inc;
wire soc_s7datacapture2_delay_slave_ce;
wire soc_s7datacapture2_serdes_m_i_delayed;
wire [7:0] soc_s7datacapture2_serdes_m_q;
wire [7:0] soc_s7datacapture2_serdes_m_d;
wire soc_s7datacapture2_serdes_s_i_delayed;
wire [7:0] soc_s7datacapture2_serdes_s_q;
wire [7:0] soc_s7datacapture2_serdes_s_d;
wire [7:0] soc_s7datacapture2_gearbox_i;
reg [9:0] soc_s7datacapture2_gearbox_o = 10'd0;
wire soc_s7datacapture2_gearbox_rst;
wire data2_cap_write_clk;
wire data2_cap_write_rst;
wire data2_cap_read_clk;
wire data2_cap_read_rst;
reg [79:0] soc_s7datacapture2_gearbox_storage = 80'd0;
reg [3:0] soc_s7datacapture2_gearbox_wrpointer = 4'd5;
reg [2:0] soc_s7datacapture2_gearbox_rdpointer = 3'd0;
wire [7:0] soc_s7datacapture2_mdata;
wire [7:0] soc_s7datacapture2_sdata;
wire soc_s7datacapture2_inc;
wire soc_s7datacapture2_dec;
wire soc_s7datacapture2_transition;
reg [7:0] soc_s7datacapture2_mdata_d = 8'd0;
reg [7:0] soc_s7datacapture2_lateness = 8'd128;
wire soc_s7datacapture2_too_late;
wire soc_s7datacapture2_too_early;
wire soc_s7datacapture2_reset_lateness;
wire soc_s7datacapture2_do_delay_rst_i;
wire soc_s7datacapture2_do_delay_rst_o;
reg soc_s7datacapture2_do_delay_rst_toggle_i = 1'd0;
wire soc_s7datacapture2_do_delay_rst_toggle_o;
reg soc_s7datacapture2_do_delay_rst_toggle_o_r = 1'd0;
wire soc_s7datacapture2_do_delay_master_inc_i;
wire soc_s7datacapture2_do_delay_master_inc_o;
reg soc_s7datacapture2_do_delay_master_inc_toggle_i = 1'd0;
wire soc_s7datacapture2_do_delay_master_inc_toggle_o;
reg soc_s7datacapture2_do_delay_master_inc_toggle_o_r = 1'd0;
wire soc_s7datacapture2_do_delay_master_dec_i;
wire soc_s7datacapture2_do_delay_master_dec_o;
reg soc_s7datacapture2_do_delay_master_dec_toggle_i = 1'd0;
wire soc_s7datacapture2_do_delay_master_dec_toggle_o;
reg soc_s7datacapture2_do_delay_master_dec_toggle_o_r = 1'd0;
wire soc_s7datacapture2_do_delay_slave_inc_i;
wire soc_s7datacapture2_do_delay_slave_inc_o;
reg soc_s7datacapture2_do_delay_slave_inc_toggle_i = 1'd0;
wire soc_s7datacapture2_do_delay_slave_inc_toggle_o;
reg soc_s7datacapture2_do_delay_slave_inc_toggle_o_r = 1'd0;
wire soc_s7datacapture2_do_delay_slave_dec_i;
wire soc_s7datacapture2_do_delay_slave_dec_o;
reg soc_s7datacapture2_do_delay_slave_dec_toggle_i = 1'd0;
wire soc_s7datacapture2_do_delay_slave_dec_toggle_o;
reg soc_s7datacapture2_do_delay_slave_dec_toggle_o_r = 1'd0;
wire soc_s7datacapture2_do_reset_lateness_i;
wire soc_s7datacapture2_do_reset_lateness_o;
reg soc_s7datacapture2_do_reset_lateness_toggle_i = 1'd0;
wire soc_s7datacapture2_do_reset_lateness_toggle_o;
reg soc_s7datacapture2_do_reset_lateness_toggle_o_r = 1'd0;
wire [9:0] soc_charsync2_raw_data;
reg soc_charsync2_synced = 1'd0;
reg [9:0] soc_charsync2_data = 10'd0;
wire soc_charsync2_char_synced_status;
wire [3:0] soc_charsync2_ctl_pos_status;
reg [9:0] soc_charsync2_raw_data1 = 10'd0;
wire [19:0] soc_charsync2_raw;
reg soc_charsync2_found_control = 1'd0;
reg [3:0] soc_charsync2_control_position = 4'd0;
reg [2:0] soc_charsync2_control_counter = 3'd0;
reg [3:0] soc_charsync2_previous_control_position = 4'd0;
reg [3:0] soc_charsync2_word_sel = 4'd0;
wire [9:0] soc_wer2_data;
wire soc_wer2_update_re;
wire soc_wer2_update_r;
reg soc_wer2_update_w = 1'd0;
reg [23:0] soc_wer2_status = 24'd0;
reg [8:0] soc_wer2_data_r = 9'd0;
reg [7:0] soc_wer2_transitions = 8'd0;
reg [3:0] soc_wer2_transition_count = 4'd0;
reg soc_wer2_is_control = 1'd0;
reg soc_wer2_is_error = 1'd0;
reg [23:0] soc_wer2_period_counter = 24'd0;
reg soc_wer2_period_done = 1'd0;
reg [23:0] soc_wer2_wer_counter = 24'd0;
reg [23:0] soc_wer2_wer_counter_r = 24'd0;
reg soc_wer2_wer_counter_r_updated = 1'd0;
reg [23:0] soc_wer2_wer_counter_sys = 24'd0;
wire soc_wer2_i;
wire soc_wer2_o;
reg soc_wer2_toggle_i = 1'd0;
wire soc_wer2_toggle_o;
reg soc_wer2_toggle_o_r = 1'd0;
wire soc_decoding2_valid_i;
wire [9:0] soc_decoding2_input;
reg soc_decoding2_valid_o = 1'd0;
reg [7:0] soc_decoding2_output_d = 8'd0;
reg [1:0] soc_decoding2_output_c = 2'd0;
reg soc_decoding2_output_de = 1'd0;
wire soc_chansync_valid_i;
reg soc_chansync_chan_synced = 1'd0;
wire soc_chansync_status;
wire soc_chansync_all_control;
wire [7:0] soc_chansync_data_in0_d;
wire [1:0] soc_chansync_data_in0_c;
wire soc_chansync_data_in0_de;
wire [7:0] soc_chansync_data_out0_d;
wire [1:0] soc_chansync_data_out0_c;
wire soc_chansync_data_out0_de;
wire [10:0] soc_chansync_syncbuffer0_din;
wire [10:0] soc_chansync_syncbuffer0_dout;
wire soc_chansync_syncbuffer0_re;
reg [2:0] soc_chansync_syncbuffer0_produce = 3'd0;
reg [2:0] soc_chansync_syncbuffer0_consume = 3'd0;
wire [2:0] soc_chansync_syncbuffer0_wrport_adr;
wire [10:0] soc_chansync_syncbuffer0_wrport_dat_r;
wire soc_chansync_syncbuffer0_wrport_we;
wire [10:0] soc_chansync_syncbuffer0_wrport_dat_w;
wire [2:0] soc_chansync_syncbuffer0_rdport_adr;
wire [10:0] soc_chansync_syncbuffer0_rdport_dat_r;
wire soc_chansync_is_control0;
wire [7:0] soc_chansync_data_in1_d;
wire [1:0] soc_chansync_data_in1_c;
wire soc_chansync_data_in1_de;
wire [7:0] soc_chansync_data_out1_d;
wire [1:0] soc_chansync_data_out1_c;
wire soc_chansync_data_out1_de;
wire [10:0] soc_chansync_syncbuffer1_din;
wire [10:0] soc_chansync_syncbuffer1_dout;
wire soc_chansync_syncbuffer1_re;
reg [2:0] soc_chansync_syncbuffer1_produce = 3'd0;
reg [2:0] soc_chansync_syncbuffer1_consume = 3'd0;
wire [2:0] soc_chansync_syncbuffer1_wrport_adr;
wire [10:0] soc_chansync_syncbuffer1_wrport_dat_r;
wire soc_chansync_syncbuffer1_wrport_we;
wire [10:0] soc_chansync_syncbuffer1_wrport_dat_w;
wire [2:0] soc_chansync_syncbuffer1_rdport_adr;
wire [10:0] soc_chansync_syncbuffer1_rdport_dat_r;
wire soc_chansync_is_control1;
wire [7:0] soc_chansync_data_in2_d;
wire [1:0] soc_chansync_data_in2_c;
wire soc_chansync_data_in2_de;
wire [7:0] soc_chansync_data_out2_d;
wire [1:0] soc_chansync_data_out2_c;
wire soc_chansync_data_out2_de;
wire [10:0] soc_chansync_syncbuffer2_din;
wire [10:0] soc_chansync_syncbuffer2_dout;
wire soc_chansync_syncbuffer2_re;
reg [2:0] soc_chansync_syncbuffer2_produce = 3'd0;
reg [2:0] soc_chansync_syncbuffer2_consume = 3'd0;
wire [2:0] soc_chansync_syncbuffer2_wrport_adr;
wire [10:0] soc_chansync_syncbuffer2_wrport_dat_r;
wire soc_chansync_syncbuffer2_wrport_we;
wire [10:0] soc_chansync_syncbuffer2_wrport_dat_w;
wire [2:0] soc_chansync_syncbuffer2_rdport_adr;
wire [10:0] soc_chansync_syncbuffer2_rdport_dat_r;
wire soc_chansync_is_control2;
wire soc_chansync_some_control;
wire soc_syncpol_valid_i;
wire [7:0] soc_syncpol_data_in0_d;
wire [1:0] soc_syncpol_data_in0_c;
wire soc_syncpol_data_in0_de;
wire [7:0] soc_syncpol_data_in1_d;
wire [1:0] soc_syncpol_data_in1_c;
wire soc_syncpol_data_in1_de;
wire [7:0] soc_syncpol_data_in2_d;
wire [1:0] soc_syncpol_data_in2_c;
wire soc_syncpol_data_in2_de;
reg soc_syncpol_valid_o = 1'd0;
wire soc_syncpol_de;
wire soc_syncpol_hsync;
wire soc_syncpol_vsync;
reg [7:0] soc_syncpol_r = 8'd0;
reg [7:0] soc_syncpol_g = 8'd0;
reg [7:0] soc_syncpol_b = 8'd0;
reg soc_syncpol_de_r = 1'd0;
reg [1:0] soc_syncpol_c_polarity = 2'd0;
reg [1:0] soc_syncpol_c_out = 2'd0;
wire soc_resdetection_valid_i;
wire soc_resdetection_vsync;
wire soc_resdetection_de;
wire [10:0] soc_resdetection_hres_status;
wire [10:0] soc_resdetection_vres_status;
reg soc_resdetection_de_r = 1'd0;
wire soc_resdetection_pn_de;
reg [10:0] soc_resdetection_hcounter = 11'd0;
reg [10:0] soc_resdetection_hcounter_st = 11'd0;
reg soc_resdetection_vsync_r = 1'd0;
wire soc_resdetection_p_vsync;
reg [10:0] soc_resdetection_vcounter = 11'd0;
reg [10:0] soc_resdetection_vcounter_st = 11'd0;
wire soc_frame_valid_i;
wire soc_frame_vsync;
wire soc_frame_de;
wire [7:0] soc_frame_r;
wire [7:0] soc_frame_g;
wire [7:0] soc_frame_b;
wire soc_frame_frame_valid;
wire soc_frame_frame_ready;
wire soc_frame_frame_first;
wire soc_frame_frame_last;
wire soc_frame_frame_payload_sof;
wire [127:0] soc_frame_frame_payload_pixels;
wire soc_frame_busy;
wire soc_frame_overflow_re;
wire soc_frame_overflow_r;
wire soc_frame_overflow_w;
reg soc_frame_de_r = 1'd0;
wire soc_frame_rgb2ycbcr_sink_valid;
wire soc_frame_rgb2ycbcr_sink_ready;
reg soc_frame_rgb2ycbcr_sink_first = 1'd0;
reg soc_frame_rgb2ycbcr_sink_last = 1'd0;
wire [7:0] soc_frame_rgb2ycbcr_sink_payload_r;
wire [7:0] soc_frame_rgb2ycbcr_sink_payload_g;
wire [7:0] soc_frame_rgb2ycbcr_sink_payload_b;
wire soc_frame_rgb2ycbcr_source_valid;
wire soc_frame_rgb2ycbcr_source_ready;
wire soc_frame_rgb2ycbcr_source_first;
wire soc_frame_rgb2ycbcr_source_last;
wire [7:0] soc_frame_rgb2ycbcr_source_payload_y;
wire [7:0] soc_frame_rgb2ycbcr_source_payload_cb;
wire [7:0] soc_frame_rgb2ycbcr_source_payload_cr;
wire [7:0] soc_frame_rgb2ycbcr_sink_r;
wire [7:0] soc_frame_rgb2ycbcr_sink_g;
wire [7:0] soc_frame_rgb2ycbcr_sink_b;
reg [7:0] soc_frame_rgb2ycbcr_source_y = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_source_cb = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_source_cr = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record0_rgb_n_r = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record0_rgb_n_g = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record0_rgb_n_b = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record1_rgb_n_r = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record1_rgb_n_g = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record1_rgb_n_b = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record2_rgb_n_r = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record2_rgb_n_g = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record2_rgb_n_b = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record3_rgb_n_r = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record3_rgb_n_g = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record3_rgb_n_b = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record4_rgb_n_r = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record4_rgb_n_g = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record4_rgb_n_b = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record5_rgb_n_r = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record5_rgb_n_g = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record5_rgb_n_b = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record6_rgb_n_r = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record6_rgb_n_g = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record6_rgb_n_b = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record7_rgb_n_r = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record7_rgb_n_g = 8'd0;
reg [7:0] soc_frame_rgb2ycbcr_record7_rgb_n_b = 8'd0;
reg signed [8:0] soc_frame_rgb2ycbcr_r_minus_g = 9'sd512;
reg signed [8:0] soc_frame_rgb2ycbcr_b_minus_g = 9'sd512;
reg signed [16:0] soc_frame_rgb2ycbcr_ca_mult_rg = 17'sd131072;
reg signed [16:0] soc_frame_rgb2ycbcr_cb_mult_bg = 17'sd131072;
reg signed [24:0] soc_frame_rgb2ycbcr_carg_plus_cbbg = 25'sd33554432;
reg signed [10:0] soc_frame_rgb2ycbcr_yraw = 11'sd2048;
reg signed [11:0] soc_frame_rgb2ycbcr_b_minus_yraw = 12'sd4096;
reg signed [11:0] soc_frame_rgb2ycbcr_r_minus_yraw = 12'sd4096;
reg signed [10:0] soc_frame_rgb2ycbcr_yraw_r0 = 11'sd2048;
reg signed [19:0] soc_frame_rgb2ycbcr_cc_mult_ryraw = 20'sd1048576;
reg signed [19:0] soc_frame_rgb2ycbcr_cd_mult_byraw = 20'sd1048576;
reg signed [10:0] soc_frame_rgb2ycbcr_yraw_r1 = 11'sd2048;
reg signed [10:0] soc_frame_rgb2ycbcr_y = 11'sd2048;
reg signed [11:0] soc_frame_rgb2ycbcr_cb = 12'sd4096;
reg signed [11:0] soc_frame_rgb2ycbcr_cr = 12'sd4096;
wire soc_frame_rgb2ycbcr_ce;
wire soc_frame_rgb2ycbcr_pipe_ce;
wire soc_frame_rgb2ycbcr_busy;
reg soc_frame_rgb2ycbcr_valid_n0 = 1'd0;
reg soc_frame_rgb2ycbcr_valid_n1 = 1'd0;
reg soc_frame_rgb2ycbcr_valid_n2 = 1'd0;
reg soc_frame_rgb2ycbcr_valid_n3 = 1'd0;
reg soc_frame_rgb2ycbcr_valid_n4 = 1'd0;
reg soc_frame_rgb2ycbcr_valid_n5 = 1'd0;
reg soc_frame_rgb2ycbcr_valid_n6 = 1'd0;
reg soc_frame_rgb2ycbcr_valid_n7 = 1'd0;
reg soc_frame_rgb2ycbcr_first_n0 = 1'd0;
reg soc_frame_rgb2ycbcr_last_n0 = 1'd0;
reg soc_frame_rgb2ycbcr_first_n1 = 1'd0;
reg soc_frame_rgb2ycbcr_last_n1 = 1'd0;
reg soc_frame_rgb2ycbcr_first_n2 = 1'd0;
reg soc_frame_rgb2ycbcr_last_n2 = 1'd0;
reg soc_frame_rgb2ycbcr_first_n3 = 1'd0;
reg soc_frame_rgb2ycbcr_last_n3 = 1'd0;
reg soc_frame_rgb2ycbcr_first_n4 = 1'd0;
reg soc_frame_rgb2ycbcr_last_n4 = 1'd0;
reg soc_frame_rgb2ycbcr_first_n5 = 1'd0;
reg soc_frame_rgb2ycbcr_last_n5 = 1'd0;
reg soc_frame_rgb2ycbcr_first_n6 = 1'd0;
reg soc_frame_rgb2ycbcr_last_n6 = 1'd0;
reg soc_frame_rgb2ycbcr_first_n7 = 1'd0;
reg soc_frame_rgb2ycbcr_last_n7 = 1'd0;
wire soc_frame_chroma_downsampler_sink_valid;
wire soc_frame_chroma_downsampler_sink_ready;
wire soc_frame_chroma_downsampler_sink_first;
wire soc_frame_chroma_downsampler_sink_last;
wire [7:0] soc_frame_chroma_downsampler_sink_payload_y;
wire [7:0] soc_frame_chroma_downsampler_sink_payload_cb;
wire [7:0] soc_frame_chroma_downsampler_sink_payload_cr;
wire soc_frame_chroma_downsampler_source_valid;
wire soc_frame_chroma_downsampler_source_ready;
wire soc_frame_chroma_downsampler_source_first;
wire soc_frame_chroma_downsampler_source_last;
wire [7:0] soc_frame_chroma_downsampler_source_payload_y;
wire [7:0] soc_frame_chroma_downsampler_source_payload_cb_cr;
wire [7:0] soc_frame_chroma_downsampler_sink_y;
wire [7:0] soc_frame_chroma_downsampler_sink_cb;
wire [7:0] soc_frame_chroma_downsampler_sink_cr;
reg [7:0] soc_frame_chroma_downsampler_source_y = 8'd0;
reg [7:0] soc_frame_chroma_downsampler_source_cb_cr = 8'd0;
wire soc_frame_chroma_downsampler_first;
reg [7:0] soc_frame_chroma_downsampler_record0_ycbcr_n_y = 8'd0;
reg [7:0] soc_frame_chroma_downsampler_record0_ycbcr_n_cb = 8'd0;
reg [7:0] soc_frame_chroma_downsampler_record0_ycbcr_n_cr = 8'd0;
reg [7:0] soc_frame_chroma_downsampler_record1_ycbcr_n_y = 8'd0;
reg [7:0] soc_frame_chroma_downsampler_record1_ycbcr_n_cb = 8'd0;
reg [7:0] soc_frame_chroma_downsampler_record1_ycbcr_n_cr = 8'd0;
reg [7:0] soc_frame_chroma_downsampler_record2_ycbcr_n_y = 8'd0;
reg [7:0] soc_frame_chroma_downsampler_record2_ycbcr_n_cb = 8'd0;
reg [7:0] soc_frame_chroma_downsampler_record2_ycbcr_n_cr = 8'd0;
reg soc_frame_chroma_downsampler_parity = 1'd0;
reg [8:0] soc_frame_chroma_downsampler_cb_sum = 9'd0;
reg [8:0] soc_frame_chroma_downsampler_cr_sum = 9'd0;
wire [7:0] soc_frame_chroma_downsampler_cb_mean;
wire [7:0] soc_frame_chroma_downsampler_cr_mean;
wire soc_frame_chroma_downsampler_ce;
wire soc_frame_chroma_downsampler_pipe_ce;
wire soc_frame_chroma_downsampler_busy;
reg soc_frame_chroma_downsampler_valid_n0 = 1'd0;
reg soc_frame_chroma_downsampler_valid_n1 = 1'd0;
reg soc_frame_chroma_downsampler_valid_n2 = 1'd0;
reg soc_frame_chroma_downsampler_first_n0 = 1'd0;
reg soc_frame_chroma_downsampler_last_n0 = 1'd0;
reg soc_frame_chroma_downsampler_first_n1 = 1'd0;
reg soc_frame_chroma_downsampler_last_n1 = 1'd0;
reg soc_frame_chroma_downsampler_first_n2 = 1'd0;
reg soc_frame_chroma_downsampler_last_n2 = 1'd0;
reg soc_frame_next_de0 = 1'd0;
reg soc_frame_next_vsync0 = 1'd0;
reg soc_frame_next_de1 = 1'd0;
reg soc_frame_next_vsync1 = 1'd0;
reg soc_frame_next_de2 = 1'd0;
reg soc_frame_next_vsync2 = 1'd0;
reg soc_frame_next_de3 = 1'd0;
reg soc_frame_next_vsync3 = 1'd0;
reg soc_frame_next_de4 = 1'd0;
reg soc_frame_next_vsync4 = 1'd0;
reg soc_frame_next_de5 = 1'd0;
reg soc_frame_next_vsync5 = 1'd0;
reg soc_frame_next_de6 = 1'd0;
reg soc_frame_next_vsync6 = 1'd0;
reg soc_frame_next_de7 = 1'd0;
reg soc_frame_next_vsync7 = 1'd0;
reg soc_frame_next_de8 = 1'd0;
reg soc_frame_next_vsync8 = 1'd0;
reg soc_frame_next_de9 = 1'd0;
reg soc_frame_next_vsync9 = 1'd0;
reg soc_frame_next_de10 = 1'd0;
reg soc_frame_next_vsync10 = 1'd0;
reg soc_frame_vsync_r = 1'd0;
wire soc_frame_new_frame;
reg [127:0] soc_frame_cur_word = 128'd0;
reg soc_frame_cur_word_valid = 1'd0;
wire [15:0] soc_frame_encoded_pixel;
reg [2:0] soc_frame_pack_counter = 3'd0;
wire soc_frame_fifo_sink_valid;
wire soc_frame_fifo_sink_ready;
reg soc_frame_fifo_sink_first = 1'd0;
reg soc_frame_fifo_sink_last = 1'd0;
reg soc_frame_fifo_sink_payload_sof = 1'd0;
wire [127:0] soc_frame_fifo_sink_payload_pixels;
wire soc_frame_fifo_source_valid;
wire soc_frame_fifo_source_ready;
wire soc_frame_fifo_source_first;
wire soc_frame_fifo_source_last;
wire soc_frame_fifo_source_payload_sof;
wire [127:0] soc_frame_fifo_source_payload_pixels;
wire soc_frame_fifo_asyncfifo_we;
wire soc_frame_fifo_asyncfifo_writable;
wire soc_frame_fifo_asyncfifo_re;
wire soc_frame_fifo_asyncfifo_readable;
wire [130:0] soc_frame_fifo_asyncfifo_din;
wire [130:0] soc_frame_fifo_asyncfifo_dout;
wire soc_frame_fifo_graycounter0_ce;
(* dont_touch = "true" *) reg [9:0] soc_frame_fifo_graycounter0_q = 10'd0;
wire [9:0] soc_frame_fifo_graycounter0_q_next;
reg [9:0] soc_frame_fifo_graycounter0_q_binary = 10'd0;
reg [9:0] soc_frame_fifo_graycounter0_q_next_binary = 10'd0;
wire soc_frame_fifo_graycounter1_ce;
(* dont_touch = "true" *) reg [9:0] soc_frame_fifo_graycounter1_q = 10'd0;
wire [9:0] soc_frame_fifo_graycounter1_q_next;
reg [9:0] soc_frame_fifo_graycounter1_q_binary = 10'd0;
reg [9:0] soc_frame_fifo_graycounter1_q_next_binary = 10'd0;
wire [9:0] soc_frame_fifo_produce_rdomain;
wire [9:0] soc_frame_fifo_consume_wdomain;
wire [8:0] soc_frame_fifo_wrport_adr;
wire [130:0] soc_frame_fifo_wrport_dat_r;
wire soc_frame_fifo_wrport_we;
wire [130:0] soc_frame_fifo_wrport_dat_w;
wire [8:0] soc_frame_fifo_rdport_adr;
wire [130:0] soc_frame_fifo_rdport_dat_r;
wire soc_frame_fifo_fifo_in_payload_sof;
wire [127:0] soc_frame_fifo_fifo_in_payload_pixels;
wire soc_frame_fifo_fifo_in_first;
wire soc_frame_fifo_fifo_in_last;
wire soc_frame_fifo_fifo_out_payload_sof;
wire [127:0] soc_frame_fifo_fifo_out_payload_pixels;
wire soc_frame_fifo_fifo_out_first;
wire soc_frame_fifo_fifo_out_last;
reg soc_frame_pix_overflow = 1'd0;
wire soc_frame_pix_overflow_reset;
wire soc_frame_sys_overflow;
wire soc_frame_overflow_reset_i;
wire soc_frame_overflow_reset_o;
reg soc_frame_overflow_reset_toggle_i = 1'd0;
wire soc_frame_overflow_reset_toggle_o;
reg soc_frame_overflow_reset_toggle_o_r = 1'd0;
wire soc_frame_overflow_reset_ack_i;
wire soc_frame_overflow_reset_ack_o;
reg soc_frame_overflow_reset_ack_toggle_i = 1'd0;
wire soc_frame_overflow_reset_ack_toggle_o;
reg soc_frame_overflow_reset_ack_toggle_o_r = 1'd0;
reg soc_frame_overflow_mask = 1'd0;
wire soc_dma_frame_valid;
reg soc_dma_frame_ready = 1'd0;
wire soc_dma_frame_first;
wire soc_dma_frame_last;
wire soc_dma_frame_payload_sof;
wire [127:0] soc_dma_frame_payload_pixels;
reg [28:0] soc_dma_frame_size_storage_full = 29'd0;
wire [24:0] soc_dma_frame_size_storage;
reg soc_dma_frame_size_re = 1'd0;
wire soc_dma_slot_array_irq;
wire [24:0] soc_dma_slot_array_address;
wire [24:0] soc_dma_slot_array_address_reached;
wire soc_dma_slot_array_address_valid;
reg soc_dma_slot_array_address_done = 1'd0;
wire soc_dma_slot_array_slot0_status;
wire soc_dma_slot_array_slot0_pending;
wire soc_dma_slot_array_slot0_trigger;
reg soc_dma_slot_array_slot0_clear = 1'd0;
wire [24:0] soc_dma_slot_array_slot0_address;
wire [24:0] soc_dma_slot_array_slot0_address_reached;
wire soc_dma_slot_array_slot0_address_valid;
wire soc_dma_slot_array_slot0_address_done;
reg [1:0] soc_dma_slot_array_slot0_status_storage_full = 2'd0;
wire [1:0] soc_dma_slot_array_slot0_status_storage;
reg soc_dma_slot_array_slot0_status_re = 1'd0;
wire soc_dma_slot_array_slot0_status_we;
wire [1:0] soc_dma_slot_array_slot0_status_dat_w;
reg [28:0] soc_dma_slot_array_slot0_address_storage_full = 29'd0;
wire [24:0] soc_dma_slot_array_slot0_address_storage;
reg soc_dma_slot_array_slot0_address_re = 1'd0;
wire soc_dma_slot_array_slot0_address_we;
wire [24:0] soc_dma_slot_array_slot0_address_dat_w;
wire soc_dma_slot_array_slot1_status;
wire soc_dma_slot_array_slot1_pending;
wire soc_dma_slot_array_slot1_trigger;
reg soc_dma_slot_array_slot1_clear = 1'd0;
wire [24:0] soc_dma_slot_array_slot1_address;
wire [24:0] soc_dma_slot_array_slot1_address_reached;
wire soc_dma_slot_array_slot1_address_valid;
wire soc_dma_slot_array_slot1_address_done;
reg [1:0] soc_dma_slot_array_slot1_status_storage_full = 2'd0;
wire [1:0] soc_dma_slot_array_slot1_status_storage;
reg soc_dma_slot_array_slot1_status_re = 1'd0;
wire soc_dma_slot_array_slot1_status_we;
wire [1:0] soc_dma_slot_array_slot1_status_dat_w;
reg [28:0] soc_dma_slot_array_slot1_address_storage_full = 29'd0;
wire [24:0] soc_dma_slot_array_slot1_address_storage;
reg soc_dma_slot_array_slot1_address_re = 1'd0;
wire soc_dma_slot_array_slot1_address_we;
wire [24:0] soc_dma_slot_array_slot1_address_dat_w;
wire soc_dma_slot_array_status_re;
wire [1:0] soc_dma_slot_array_status_r;
reg [1:0] soc_dma_slot_array_status_w = 2'd0;
wire soc_dma_slot_array_pending_re;
wire [1:0] soc_dma_slot_array_pending_r;
reg [1:0] soc_dma_slot_array_pending_w = 2'd0;
reg [1:0] soc_dma_slot_array_storage_full = 2'd0;
wire [1:0] soc_dma_slot_array_storage;
reg soc_dma_slot_array_re = 1'd0;
wire soc_dma_slot_array_change_slot;
reg soc_dma_slot_array_current_slot = 1'd0;
reg soc_dma_reset_words = 1'd0;
reg soc_dma_count_word = 1'd0;
wire soc_dma_last_word;
reg [24:0] soc_dma_current_address = 25'd0;
reg [24:0] soc_dma_mwords_remaining = 25'd0;
wire [127:0] soc_dma_memory_word;
reg soc_dma_sink_sink_valid = 1'd0;
wire soc_dma_sink_sink_ready;
wire [24:0] soc_dma_sink_sink_payload_address;
wire [127:0] soc_dma_sink_sink_payload_data;
wire soc_dma_fifo_sink_valid;
wire soc_dma_fifo_sink_ready;
reg soc_dma_fifo_sink_first = 1'd0;
reg soc_dma_fifo_sink_last = 1'd0;
wire [127:0] soc_dma_fifo_sink_payload_data;
wire soc_dma_fifo_source_valid;
wire soc_dma_fifo_source_ready;
wire soc_dma_fifo_source_first;
wire soc_dma_fifo_source_last;
wire [127:0] soc_dma_fifo_source_payload_data;
wire soc_dma_fifo_syncfifo_we;
wire soc_dma_fifo_syncfifo_writable;
wire soc_dma_fifo_syncfifo_re;
wire soc_dma_fifo_syncfifo_readable;
wire [129:0] soc_dma_fifo_syncfifo_din;
wire [129:0] soc_dma_fifo_syncfifo_dout;
reg [4:0] soc_dma_fifo_level = 5'd0;
reg soc_dma_fifo_replace = 1'd0;
reg [3:0] soc_dma_fifo_produce = 4'd0;
reg [3:0] soc_dma_fifo_consume = 4'd0;
reg [3:0] soc_dma_fifo_wrport_adr = 4'd0;
wire [129:0] soc_dma_fifo_wrport_dat_r;
wire soc_dma_fifo_wrport_we;
wire [129:0] soc_dma_fifo_wrport_dat_w;
wire soc_dma_fifo_do_read;
wire [3:0] soc_dma_fifo_rdport_adr;
wire [129:0] soc_dma_fifo_rdport_dat_r;
wire [127:0] soc_dma_fifo_fifo_in_payload_data;
wire soc_dma_fifo_fifo_in_first;
wire soc_dma_fifo_fifo_in_last;
wire [127:0] soc_dma_fifo_fifo_out_payload_data;
wire soc_dma_fifo_fifo_out_first;
wire soc_dma_fifo_fifo_out_last;
wire soc_hdmi_in0_freq_clk0;
wire [31:0] soc_hdmi_in0_freq_status;
wire fmeter_clk;
wire soc_hdmi_in0_freq_period_done;
reg [31:0] soc_hdmi_in0_freq_period_counter = 32'd0;
wire soc_hdmi_in0_freq_ce;
reg [5:0] soc_hdmi_in0_freq_q = 6'd0;
wire [5:0] soc_hdmi_in0_freq_q_next;
reg [5:0] soc_hdmi_in0_freq_q_binary = 6'd0;
reg [5:0] soc_hdmi_in0_freq_q_next_binary = 6'd0;
wire [5:0] soc_hdmi_in0_freq_gray_decoder_i;
reg [5:0] soc_hdmi_in0_freq_gray_decoder_o = 6'd0;
reg [5:0] soc_hdmi_in0_freq_gray_decoder_o_comb = 6'd0;
wire soc_hdmi_in0_freq_sampler_latch;
wire [5:0] soc_hdmi_in0_freq_sampler_i;
reg [31:0] soc_hdmi_in0_freq_sampler_o = 32'd0;
wire [5:0] soc_hdmi_in0_freq_sampler_inc;
reg [31:0] soc_hdmi_in0_freq_sampler_counter = 32'd0;
reg [5:0] soc_hdmi_in0_freq_sampler_i_d = 6'd0;
wire soc_hdmi_out0_dram_port_cmd_valid;
wire soc_hdmi_out0_dram_port_cmd_ready;
wire soc_hdmi_out0_dram_port_cmd_first;
wire soc_hdmi_out0_dram_port_cmd_last;
wire soc_hdmi_out0_dram_port_cmd_payload_we;
wire [24:0] soc_hdmi_out0_dram_port_cmd_payload_adr;
wire soc_hdmi_out0_dram_port_wdata_ready;
reg [127:0] soc_hdmi_out0_dram_port_wdata_payload_data = 128'd0;
reg [15:0] soc_hdmi_out0_dram_port_wdata_payload_we = 16'd0;
wire soc_hdmi_out0_dram_port_rdata_valid;
wire soc_hdmi_out0_dram_port_rdata_ready;
reg soc_hdmi_out0_dram_port_rdata_first = 1'd0;
reg soc_hdmi_out0_dram_port_rdata_last = 1'd0;
wire [127:0] soc_hdmi_out0_dram_port_rdata_payload_data;
reg soc_hdmi_out0_dram_port_litedramport0_cmd_valid = 1'd0;
wire soc_hdmi_out0_dram_port_litedramport0_cmd_ready;
reg soc_hdmi_out0_dram_port_litedramport0_cmd_first = 1'd0;
reg soc_hdmi_out0_dram_port_litedramport0_cmd_last = 1'd0;
reg soc_hdmi_out0_dram_port_litedramport0_cmd_payload_we = 1'd0;
reg [24:0] soc_hdmi_out0_dram_port_litedramport0_cmd_payload_adr = 25'd0;
wire soc_hdmi_out0_dram_port_litedramport0_rdata_valid;
wire soc_hdmi_out0_dram_port_litedramport0_rdata_ready;
wire soc_hdmi_out0_dram_port_litedramport0_rdata_first;
wire soc_hdmi_out0_dram_port_litedramport0_rdata_last;
wire [127:0] soc_hdmi_out0_dram_port_litedramport0_rdata_payload_data;
wire soc_hdmi_out0_dram_port_cmd_fifo_sink_valid;
wire soc_hdmi_out0_dram_port_cmd_fifo_sink_ready;
wire soc_hdmi_out0_dram_port_cmd_fifo_sink_first;
wire soc_hdmi_out0_dram_port_cmd_fifo_sink_last;
wire soc_hdmi_out0_dram_port_cmd_fifo_sink_payload_we;
wire [24:0] soc_hdmi_out0_dram_port_cmd_fifo_sink_payload_adr;
wire soc_hdmi_out0_dram_port_cmd_fifo_source_valid;
wire soc_hdmi_out0_dram_port_cmd_fifo_source_ready;
wire soc_hdmi_out0_dram_port_cmd_fifo_source_first;
wire soc_hdmi_out0_dram_port_cmd_fifo_source_last;
wire soc_hdmi_out0_dram_port_cmd_fifo_source_payload_we;
wire [24:0] soc_hdmi_out0_dram_port_cmd_fifo_source_payload_adr;
wire soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_we;
wire soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_writable;
wire soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_re;
wire soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_readable;
wire [27:0] soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_din;
wire [27:0] soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_dout;
wire soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_ce;
(* dont_touch = "true" *) reg [2:0] soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q = 3'd0;
wire [2:0] soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next;
reg [2:0] soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_binary = 3'd0;
reg [2:0] soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next_binary = 3'd0;
wire soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_ce;
(* dont_touch = "true" *) reg [2:0] soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q = 3'd0;
wire [2:0] soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next;
reg [2:0] soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_binary = 3'd0;
reg [2:0] soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary = 3'd0;
wire [2:0] soc_hdmi_out0_dram_port_cmd_fifo_produce_rdomain;
wire [2:0] soc_hdmi_out0_dram_port_cmd_fifo_consume_wdomain;
wire [1:0] soc_hdmi_out0_dram_port_cmd_fifo_wrport_adr;
wire [27:0] soc_hdmi_out0_dram_port_cmd_fifo_wrport_dat_r;
wire soc_hdmi_out0_dram_port_cmd_fifo_wrport_we;
wire [27:0] soc_hdmi_out0_dram_port_cmd_fifo_wrport_dat_w;
wire [1:0] soc_hdmi_out0_dram_port_cmd_fifo_rdport_adr;
wire [27:0] soc_hdmi_out0_dram_port_cmd_fifo_rdport_dat_r;
wire soc_hdmi_out0_dram_port_cmd_fifo_fifo_in_payload_we;
wire [24:0] soc_hdmi_out0_dram_port_cmd_fifo_fifo_in_payload_adr;
wire soc_hdmi_out0_dram_port_cmd_fifo_fifo_in_first;
wire soc_hdmi_out0_dram_port_cmd_fifo_fifo_in_last;
wire soc_hdmi_out0_dram_port_cmd_fifo_fifo_out_payload_we;
wire [24:0] soc_hdmi_out0_dram_port_cmd_fifo_fifo_out_payload_adr;
wire soc_hdmi_out0_dram_port_cmd_fifo_fifo_out_first;
wire soc_hdmi_out0_dram_port_cmd_fifo_fifo_out_last;
wire soc_hdmi_out0_dram_port_rdata_fifo_sink_valid;
wire soc_hdmi_out0_dram_port_rdata_fifo_sink_ready;
wire soc_hdmi_out0_dram_port_rdata_fifo_sink_first;
wire soc_hdmi_out0_dram_port_rdata_fifo_sink_last;
wire [127:0] soc_hdmi_out0_dram_port_rdata_fifo_sink_payload_data;
wire soc_hdmi_out0_dram_port_rdata_fifo_source_valid;
wire soc_hdmi_out0_dram_port_rdata_fifo_source_ready;
wire soc_hdmi_out0_dram_port_rdata_fifo_source_first;
wire soc_hdmi_out0_dram_port_rdata_fifo_source_last;
wire [127:0] soc_hdmi_out0_dram_port_rdata_fifo_source_payload_data;
wire soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_we;
wire soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_writable;
wire soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_re;
wire soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_readable;
wire [129:0] soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_din;
wire [129:0] soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_dout;
wire soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_ce;
(* dont_touch = "true" *) reg [4:0] soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q = 5'd0;
wire [4:0] soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next;
reg [4:0] soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_binary = 5'd0;
reg [4:0] soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next_binary = 5'd0;
wire soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_ce;
(* dont_touch = "true" *) reg [4:0] soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q = 5'd0;
wire [4:0] soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next;
reg [4:0] soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_binary = 5'd0;
reg [4:0] soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary = 5'd0;
wire [4:0] soc_hdmi_out0_dram_port_rdata_fifo_produce_rdomain;
wire [4:0] soc_hdmi_out0_dram_port_rdata_fifo_consume_wdomain;
wire [3:0] soc_hdmi_out0_dram_port_rdata_fifo_wrport_adr;
wire [129:0] soc_hdmi_out0_dram_port_rdata_fifo_wrport_dat_r;
wire soc_hdmi_out0_dram_port_rdata_fifo_wrport_we;
wire [129:0] soc_hdmi_out0_dram_port_rdata_fifo_wrport_dat_w;
wire [3:0] soc_hdmi_out0_dram_port_rdata_fifo_rdport_adr;
wire [129:0] soc_hdmi_out0_dram_port_rdata_fifo_rdport_dat_r;
wire [127:0] soc_hdmi_out0_dram_port_rdata_fifo_fifo_in_payload_data;
wire soc_hdmi_out0_dram_port_rdata_fifo_fifo_in_first;
wire soc_hdmi_out0_dram_port_rdata_fifo_fifo_in_last;
wire [127:0] soc_hdmi_out0_dram_port_rdata_fifo_fifo_out_payload_data;
wire soc_hdmi_out0_dram_port_rdata_fifo_fifo_out_first;
wire soc_hdmi_out0_dram_port_rdata_fifo_fifo_out_last;
wire soc_hdmi_out0_dram_port_litedramport1_cmd_valid;
reg soc_hdmi_out0_dram_port_litedramport1_cmd_ready = 1'd0;
wire soc_hdmi_out0_dram_port_litedramport1_cmd_payload_we;
wire [27:0] soc_hdmi_out0_dram_port_litedramport1_cmd_payload_adr;
reg soc_hdmi_out0_dram_port_litedramport1_rdata_valid = 1'd0;
wire soc_hdmi_out0_dram_port_litedramport1_rdata_ready;
reg soc_hdmi_out0_dram_port_litedramport1_rdata_first = 1'd0;
reg soc_hdmi_out0_dram_port_litedramport1_rdata_last = 1'd0;
reg [15:0] soc_hdmi_out0_dram_port_litedramport1_rdata_payload_data = 16'd0;
reg soc_hdmi_out0_dram_port_litedramport1_flush = 1'd0;
reg soc_hdmi_out0_dram_port_cmd_buffer_sink_valid = 1'd0;
wire soc_hdmi_out0_dram_port_cmd_buffer_sink_ready;
reg soc_hdmi_out0_dram_port_cmd_buffer_sink_first = 1'd0;
reg soc_hdmi_out0_dram_port_cmd_buffer_sink_last = 1'd0;
reg [7:0] soc_hdmi_out0_dram_port_cmd_buffer_sink_payload_sel = 8'd0;
wire soc_hdmi_out0_dram_port_cmd_buffer_source_valid;
wire soc_hdmi_out0_dram_port_cmd_buffer_source_ready;
wire soc_hdmi_out0_dram_port_cmd_buffer_source_first;
wire soc_hdmi_out0_dram_port_cmd_buffer_source_last;
wire [7:0] soc_hdmi_out0_dram_port_cmd_buffer_source_payload_sel;
wire soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_we;
wire soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_writable;
wire soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_re;
wire soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_readable;
wire [9:0] soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_din;
wire [9:0] soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_dout;
reg [2:0] soc_hdmi_out0_dram_port_cmd_buffer_level = 3'd0;
reg soc_hdmi_out0_dram_port_cmd_buffer_replace = 1'd0;
reg [1:0] soc_hdmi_out0_dram_port_cmd_buffer_produce = 2'd0;
reg [1:0] soc_hdmi_out0_dram_port_cmd_buffer_consume = 2'd0;
reg [1:0] soc_hdmi_out0_dram_port_cmd_buffer_wrport_adr = 2'd0;
wire [9:0] soc_hdmi_out0_dram_port_cmd_buffer_wrport_dat_r;
wire soc_hdmi_out0_dram_port_cmd_buffer_wrport_we;
wire [9:0] soc_hdmi_out0_dram_port_cmd_buffer_wrport_dat_w;
wire soc_hdmi_out0_dram_port_cmd_buffer_do_read;
wire [1:0] soc_hdmi_out0_dram_port_cmd_buffer_rdport_adr;
wire [9:0] soc_hdmi_out0_dram_port_cmd_buffer_rdport_dat_r;
wire [7:0] soc_hdmi_out0_dram_port_cmd_buffer_fifo_in_payload_sel;
wire soc_hdmi_out0_dram_port_cmd_buffer_fifo_in_first;
wire soc_hdmi_out0_dram_port_cmd_buffer_fifo_in_last;
wire [7:0] soc_hdmi_out0_dram_port_cmd_buffer_fifo_out_payload_sel;
wire soc_hdmi_out0_dram_port_cmd_buffer_fifo_out_first;
wire soc_hdmi_out0_dram_port_cmd_buffer_fifo_out_last;
reg [2:0] soc_hdmi_out0_dram_port_counter = 3'd0;
reg soc_hdmi_out0_dram_port_counter_ce = 1'd0;
wire soc_hdmi_out0_dram_port_rdata_buffer_sink_valid;
wire soc_hdmi_out0_dram_port_rdata_buffer_sink_ready;
wire soc_hdmi_out0_dram_port_rdata_buffer_sink_first;
wire soc_hdmi_out0_dram_port_rdata_buffer_sink_last;
wire [127:0] soc_hdmi_out0_dram_port_rdata_buffer_sink_payload_data;
wire soc_hdmi_out0_dram_port_rdata_buffer_source_valid;
wire soc_hdmi_out0_dram_port_rdata_buffer_source_ready;
wire soc_hdmi_out0_dram_port_rdata_buffer_source_first;
wire soc_hdmi_out0_dram_port_rdata_buffer_source_last;
reg [127:0] soc_hdmi_out0_dram_port_rdata_buffer_source_payload_data = 128'd0;
wire soc_hdmi_out0_dram_port_rdata_buffer_pipe_ce;
wire soc_hdmi_out0_dram_port_rdata_buffer_busy;
reg soc_hdmi_out0_dram_port_rdata_buffer_valid_n = 1'd0;
reg soc_hdmi_out0_dram_port_rdata_buffer_first_n = 1'd0;
reg soc_hdmi_out0_dram_port_rdata_buffer_last_n = 1'd0;
wire soc_hdmi_out0_dram_port_rdata_converter_sink_valid;
wire soc_hdmi_out0_dram_port_rdata_converter_sink_ready;
wire soc_hdmi_out0_dram_port_rdata_converter_sink_first;
wire soc_hdmi_out0_dram_port_rdata_converter_sink_last;
wire [127:0] soc_hdmi_out0_dram_port_rdata_converter_sink_payload_data;
wire soc_hdmi_out0_dram_port_rdata_converter_source_valid;
reg soc_hdmi_out0_dram_port_rdata_converter_source_ready = 1'd0;
wire soc_hdmi_out0_dram_port_rdata_converter_source_first;
wire soc_hdmi_out0_dram_port_rdata_converter_source_last;
wire [15:0] soc_hdmi_out0_dram_port_rdata_converter_source_payload_data;
wire soc_hdmi_out0_dram_port_rdata_converter_converter_sink_valid;
wire soc_hdmi_out0_dram_port_rdata_converter_converter_sink_ready;
wire soc_hdmi_out0_dram_port_rdata_converter_converter_sink_first;
wire soc_hdmi_out0_dram_port_rdata_converter_converter_sink_last;
reg [127:0] soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data = 128'd0;
wire soc_hdmi_out0_dram_port_rdata_converter_converter_source_valid;
wire soc_hdmi_out0_dram_port_rdata_converter_converter_source_ready;
wire soc_hdmi_out0_dram_port_rdata_converter_converter_source_first;
wire soc_hdmi_out0_dram_port_rdata_converter_converter_source_last;
reg [15:0] soc_hdmi_out0_dram_port_rdata_converter_converter_source_payload_data = 16'd0;
wire soc_hdmi_out0_dram_port_rdata_converter_converter_source_payload_valid_token_count;
reg [2:0] soc_hdmi_out0_dram_port_rdata_converter_converter_mux = 3'd0;
wire soc_hdmi_out0_dram_port_rdata_converter_converter_first;
wire soc_hdmi_out0_dram_port_rdata_converter_converter_last;
wire soc_hdmi_out0_dram_port_rdata_converter_source_source_valid;
wire soc_hdmi_out0_dram_port_rdata_converter_source_source_ready;
wire soc_hdmi_out0_dram_port_rdata_converter_source_source_first;
wire soc_hdmi_out0_dram_port_rdata_converter_source_source_last;
wire [15:0] soc_hdmi_out0_dram_port_rdata_converter_source_source_payload_data;
reg [7:0] soc_hdmi_out0_dram_port_rdata_chunk = 8'd1;
wire soc_hdmi_out0_dram_port_rdata_chunk_valid;
wire soc_hdmi_out0_core_source_source_valid;
wire soc_hdmi_out0_core_source_source_ready;
wire [15:0] soc_hdmi_out0_core_source_source_payload_data;
wire soc_hdmi_out0_core_source_source_param_hsync;
wire soc_hdmi_out0_core_source_source_param_vsync;
wire soc_hdmi_out0_core_source_source_param_de;
reg soc_hdmi_out0_core_underflow_enable_storage_full = 1'd0;
wire soc_hdmi_out0_core_underflow_enable_storage;
reg soc_hdmi_out0_core_underflow_enable_re = 1'd0;
wire soc_hdmi_out0_core_underflow_update_underflow_update_re;
wire soc_hdmi_out0_core_underflow_update_underflow_update_r;
reg soc_hdmi_out0_core_underflow_update_underflow_update_w = 1'd0;
reg [31:0] soc_hdmi_out0_core_underflow_counter_status = 32'd0;
wire soc_hdmi_out0_core_initiator_source_source_valid;
wire soc_hdmi_out0_core_initiator_source_source_ready;
wire soc_hdmi_out0_core_initiator_source_source_first;
wire soc_hdmi_out0_core_initiator_source_source_last;
wire [11:0] soc_hdmi_out0_core_initiator_source_source_payload_hres;
wire [11:0] soc_hdmi_out0_core_initiator_source_source_payload_hsync_start;
wire [11:0] soc_hdmi_out0_core_initiator_source_source_payload_hsync_end;
wire [11:0] soc_hdmi_out0_core_initiator_source_source_payload_hscan;
wire [11:0] soc_hdmi_out0_core_initiator_source_source_payload_vres;
wire [11:0] soc_hdmi_out0_core_initiator_source_source_payload_vsync_start;
wire [11:0] soc_hdmi_out0_core_initiator_source_source_payload_vsync_end;
wire [11:0] soc_hdmi_out0_core_initiator_source_source_payload_vscan;
wire [31:0] soc_hdmi_out0_core_initiator_source_source_payload_base;
wire [31:0] soc_hdmi_out0_core_initiator_source_source_payload_length;
wire soc_hdmi_out0_core_initiator_cdc_sink_valid;
wire soc_hdmi_out0_core_initiator_cdc_sink_ready;
reg soc_hdmi_out0_core_initiator_cdc_sink_first = 1'd0;
reg soc_hdmi_out0_core_initiator_cdc_sink_last = 1'd0;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_sink_payload_hres;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_sink_payload_hsync_start;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_sink_payload_hsync_end;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_sink_payload_hscan;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_sink_payload_vres;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_sink_payload_vsync_start;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_sink_payload_vsync_end;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_sink_payload_vscan;
wire [31:0] soc_hdmi_out0_core_initiator_cdc_sink_payload_base;
wire [31:0] soc_hdmi_out0_core_initiator_cdc_sink_payload_length;
wire soc_hdmi_out0_core_initiator_cdc_source_valid;
wire soc_hdmi_out0_core_initiator_cdc_source_ready;
wire soc_hdmi_out0_core_initiator_cdc_source_first;
wire soc_hdmi_out0_core_initiator_cdc_source_last;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_source_payload_hres;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_source_payload_hsync_start;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_source_payload_hsync_end;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_source_payload_hscan;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_source_payload_vres;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_source_payload_vsync_start;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_source_payload_vsync_end;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_source_payload_vscan;
wire [31:0] soc_hdmi_out0_core_initiator_cdc_source_payload_base;
wire [31:0] soc_hdmi_out0_core_initiator_cdc_source_payload_length;
wire soc_hdmi_out0_core_initiator_cdc_asyncfifo_we;
wire soc_hdmi_out0_core_initiator_cdc_asyncfifo_writable;
wire soc_hdmi_out0_core_initiator_cdc_asyncfifo_re;
wire soc_hdmi_out0_core_initiator_cdc_asyncfifo_readable;
wire [161:0] soc_hdmi_out0_core_initiator_cdc_asyncfifo_din;
wire [161:0] soc_hdmi_out0_core_initiator_cdc_asyncfifo_dout;
wire soc_hdmi_out0_core_initiator_cdc_graycounter0_ce;
(* dont_touch = "true" *) reg [1:0] soc_hdmi_out0_core_initiator_cdc_graycounter0_q = 2'd0;
wire [1:0] soc_hdmi_out0_core_initiator_cdc_graycounter0_q_next;
reg [1:0] soc_hdmi_out0_core_initiator_cdc_graycounter0_q_binary = 2'd0;
reg [1:0] soc_hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary = 2'd0;
wire soc_hdmi_out0_core_initiator_cdc_graycounter1_ce;
(* dont_touch = "true" *) reg [1:0] soc_hdmi_out0_core_initiator_cdc_graycounter1_q = 2'd0;
wire [1:0] soc_hdmi_out0_core_initiator_cdc_graycounter1_q_next;
reg [1:0] soc_hdmi_out0_core_initiator_cdc_graycounter1_q_binary = 2'd0;
reg [1:0] soc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary = 2'd0;
wire [1:0] soc_hdmi_out0_core_initiator_cdc_produce_rdomain;
wire [1:0] soc_hdmi_out0_core_initiator_cdc_consume_wdomain;
wire soc_hdmi_out0_core_initiator_cdc_wrport_adr;
wire [161:0] soc_hdmi_out0_core_initiator_cdc_wrport_dat_r;
wire soc_hdmi_out0_core_initiator_cdc_wrport_we;
wire [161:0] soc_hdmi_out0_core_initiator_cdc_wrport_dat_w;
wire soc_hdmi_out0_core_initiator_cdc_rdport_adr;
wire [161:0] soc_hdmi_out0_core_initiator_cdc_rdport_dat_r;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hres;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_start;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_end;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hscan;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vres;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_start;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_end;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vscan;
wire [31:0] soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_base;
wire [31:0] soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_length;
wire soc_hdmi_out0_core_initiator_cdc_fifo_in_first;
wire soc_hdmi_out0_core_initiator_cdc_fifo_in_last;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hres;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_start;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_end;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hscan;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vres;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_start;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_end;
wire [11:0] soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vscan;
wire [31:0] soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_base;
wire [31:0] soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_length;
wire soc_hdmi_out0_core_initiator_cdc_fifo_out_first;
wire soc_hdmi_out0_core_initiator_cdc_fifo_out_last;
reg soc_hdmi_out0_core_initiator_enable_storage_full = 1'd0;
wire soc_hdmi_out0_core_initiator_enable_storage;
reg soc_hdmi_out0_core_initiator_enable_re = 1'd0;
reg [11:0] soc_hdmi_out0_core_initiator_csrstorage0_storage_full = 12'd0;
wire [11:0] soc_hdmi_out0_core_initiator_csrstorage0_storage;
reg soc_hdmi_out0_core_initiator_csrstorage0_re = 1'd0;
reg [11:0] soc_hdmi_out0_core_initiator_csrstorage1_storage_full = 12'd0;
wire [11:0] soc_hdmi_out0_core_initiator_csrstorage1_storage;
reg soc_hdmi_out0_core_initiator_csrstorage1_re = 1'd0;
reg [11:0] soc_hdmi_out0_core_initiator_csrstorage2_storage_full = 12'd0;
wire [11:0] soc_hdmi_out0_core_initiator_csrstorage2_storage;
reg soc_hdmi_out0_core_initiator_csrstorage2_re = 1'd0;
reg [11:0] soc_hdmi_out0_core_initiator_csrstorage3_storage_full = 12'd0;
wire [11:0] soc_hdmi_out0_core_initiator_csrstorage3_storage;
reg soc_hdmi_out0_core_initiator_csrstorage3_re = 1'd0;
reg [11:0] soc_hdmi_out0_core_initiator_csrstorage4_storage_full = 12'd0;
wire [11:0] soc_hdmi_out0_core_initiator_csrstorage4_storage;
reg soc_hdmi_out0_core_initiator_csrstorage4_re = 1'd0;
reg [11:0] soc_hdmi_out0_core_initiator_csrstorage5_storage_full = 12'd0;
wire [11:0] soc_hdmi_out0_core_initiator_csrstorage5_storage;
reg soc_hdmi_out0_core_initiator_csrstorage5_re = 1'd0;
reg [11:0] soc_hdmi_out0_core_initiator_csrstorage6_storage_full = 12'd0;
wire [11:0] soc_hdmi_out0_core_initiator_csrstorage6_storage;
reg soc_hdmi_out0_core_initiator_csrstorage6_re = 1'd0;
reg [11:0] soc_hdmi_out0_core_initiator_csrstorage7_storage_full = 12'd0;
wire [11:0] soc_hdmi_out0_core_initiator_csrstorage7_storage;
reg soc_hdmi_out0_core_initiator_csrstorage7_re = 1'd0;
reg [31:0] soc_hdmi_out0_core_initiator_csrstorage8_storage_full = 32'd0;
wire [31:0] soc_hdmi_out0_core_initiator_csrstorage8_storage;
reg soc_hdmi_out0_core_initiator_csrstorage8_re = 1'd0;
reg [31:0] soc_hdmi_out0_core_initiator_csrstorage9_storage_full = 32'd0;
wire [31:0] soc_hdmi_out0_core_initiator_csrstorage9_storage;
reg soc_hdmi_out0_core_initiator_csrstorage9_re = 1'd0;
wire soc_hdmi_out0_core_timinggenerator_sink_valid;
wire soc_hdmi_out0_core_timinggenerator_sink_ready;
wire [11:0] soc_hdmi_out0_core_timinggenerator_sink_payload_hres;
wire [11:0] soc_hdmi_out0_core_timinggenerator_sink_payload_hsync_start;
wire [11:0] soc_hdmi_out0_core_timinggenerator_sink_payload_hsync_end;
wire [11:0] soc_hdmi_out0_core_timinggenerator_sink_payload_hscan;
wire [11:0] soc_hdmi_out0_core_timinggenerator_sink_payload_vres;
wire [11:0] soc_hdmi_out0_core_timinggenerator_sink_payload_vsync_start;
wire [11:0] soc_hdmi_out0_core_timinggenerator_sink_payload_vsync_end;
wire [11:0] soc_hdmi_out0_core_timinggenerator_sink_payload_vscan;
reg soc_hdmi_out0_core_timinggenerator_source_valid = 1'd0;
reg soc_hdmi_out0_core_timinggenerator_source_ready = 1'd0;
reg soc_hdmi_out0_core_timinggenerator_source_last = 1'd0;
reg soc_hdmi_out0_core_timinggenerator_source_payload_hsync = 1'd0;
reg soc_hdmi_out0_core_timinggenerator_source_payload_vsync = 1'd0;
reg soc_hdmi_out0_core_timinggenerator_source_payload_de = 1'd0;
reg soc_hdmi_out0_core_timinggenerator_hactive = 1'd0;
reg soc_hdmi_out0_core_timinggenerator_vactive = 1'd0;
reg soc_hdmi_out0_core_timinggenerator_active = 1'd0;
reg [11:0] soc_hdmi_out0_core_timinggenerator_hcounter = 12'd0;
reg [11:0] soc_hdmi_out0_core_timinggenerator_vcounter = 12'd0;
wire soc_hdmi_out0_core_dmareader_sink_valid;
reg soc_hdmi_out0_core_dmareader_sink_ready = 1'd0;
wire [31:0] soc_hdmi_out0_core_dmareader_sink_payload_base;
wire [31:0] soc_hdmi_out0_core_dmareader_sink_payload_length;
wire soc_hdmi_out0_core_dmareader_source_valid;
reg soc_hdmi_out0_core_dmareader_source_ready = 1'd0;
wire soc_hdmi_out0_core_dmareader_source_first;
wire soc_hdmi_out0_core_dmareader_source_last;
wire [15:0] soc_hdmi_out0_core_dmareader_source_payload_data;
reg soc_hdmi_out0_core_dmareader_sink_sink_valid = 1'd0;
wire soc_hdmi_out0_core_dmareader_sink_sink_ready;
wire [27:0] soc_hdmi_out0_core_dmareader_sink_sink_payload_address;
wire soc_hdmi_out0_core_dmareader_source_source_valid;
wire soc_hdmi_out0_core_dmareader_source_source_ready;
wire soc_hdmi_out0_core_dmareader_source_source_first;
wire soc_hdmi_out0_core_dmareader_source_source_last;
wire [15:0] soc_hdmi_out0_core_dmareader_source_source_payload_data;
wire soc_hdmi_out0_core_dmareader_request_enable;
wire soc_hdmi_out0_core_dmareader_request_issued;
wire soc_hdmi_out0_core_dmareader_data_dequeued;
reg [12:0] soc_hdmi_out0_core_dmareader_rsv_level = 13'd0;
wire soc_hdmi_out0_core_dmareader_fifo_sink_valid;
wire soc_hdmi_out0_core_dmareader_fifo_sink_ready;
wire soc_hdmi_out0_core_dmareader_fifo_sink_first;
wire soc_hdmi_out0_core_dmareader_fifo_sink_last;
wire [15:0] soc_hdmi_out0_core_dmareader_fifo_sink_payload_data;
wire soc_hdmi_out0_core_dmareader_fifo_source_valid;
wire soc_hdmi_out0_core_dmareader_fifo_source_ready;
wire soc_hdmi_out0_core_dmareader_fifo_source_first;
wire soc_hdmi_out0_core_dmareader_fifo_source_last;
wire [15:0] soc_hdmi_out0_core_dmareader_fifo_source_payload_data;
wire soc_hdmi_out0_core_dmareader_fifo_re;
reg soc_hdmi_out0_core_dmareader_fifo_readable = 1'd0;
wire soc_hdmi_out0_core_dmareader_fifo_syncfifo_we;
wire soc_hdmi_out0_core_dmareader_fifo_syncfifo_writable;
wire soc_hdmi_out0_core_dmareader_fifo_syncfifo_re;
wire soc_hdmi_out0_core_dmareader_fifo_syncfifo_readable;
wire [17:0] soc_hdmi_out0_core_dmareader_fifo_syncfifo_din;
wire [17:0] soc_hdmi_out0_core_dmareader_fifo_syncfifo_dout;
reg [12:0] soc_hdmi_out0_core_dmareader_fifo_level0 = 13'd0;
reg soc_hdmi_out0_core_dmareader_fifo_replace = 1'd0;
reg [11:0] soc_hdmi_out0_core_dmareader_fifo_produce = 12'd0;
reg [11:0] soc_hdmi_out0_core_dmareader_fifo_consume = 12'd0;
reg [11:0] soc_hdmi_out0_core_dmareader_fifo_wrport_adr = 12'd0;
wire [17:0] soc_hdmi_out0_core_dmareader_fifo_wrport_dat_r;
wire soc_hdmi_out0_core_dmareader_fifo_wrport_we;
wire [17:0] soc_hdmi_out0_core_dmareader_fifo_wrport_dat_w;
wire soc_hdmi_out0_core_dmareader_fifo_do_read;
wire [11:0] soc_hdmi_out0_core_dmareader_fifo_rdport_adr;
wire [17:0] soc_hdmi_out0_core_dmareader_fifo_rdport_dat_r;
wire soc_hdmi_out0_core_dmareader_fifo_rdport_re;
wire [12:0] soc_hdmi_out0_core_dmareader_fifo_level1;
wire [15:0] soc_hdmi_out0_core_dmareader_fifo_fifo_in_payload_data;
wire soc_hdmi_out0_core_dmareader_fifo_fifo_in_first;
wire soc_hdmi_out0_core_dmareader_fifo_fifo_in_last;
wire [15:0] soc_hdmi_out0_core_dmareader_fifo_fifo_out_payload_data;
wire soc_hdmi_out0_core_dmareader_fifo_fifo_out_first;
wire soc_hdmi_out0_core_dmareader_fifo_fifo_out_last;
wire [27:0] soc_hdmi_out0_core_dmareader_base;
wire [27:0] soc_hdmi_out0_core_dmareader_length;
reg [27:0] soc_hdmi_out0_core_dmareader_offset = 28'd0;
wire soc_hdmi_out0_core_underflow_enable;
wire soc_hdmi_out0_core_underflow_update;
reg [31:0] soc_hdmi_out0_core_underflow_counter = 32'd0;
wire soc_hdmi_out0_core_i;
wire soc_hdmi_out0_core_o;
reg soc_hdmi_out0_core_toggle_i = 1'd0;
wire soc_hdmi_out0_core_toggle_o;
reg soc_hdmi_out0_core_toggle_o_r = 1'd0;
wire soc_hdmi_out0_driver_sink_sink_valid;
wire soc_hdmi_out0_driver_sink_sink_ready;
wire soc_hdmi_out0_driver_sink_sink_first;
wire soc_hdmi_out0_driver_sink_sink_last;
wire [7:0] soc_hdmi_out0_driver_sink_sink_payload_r;
wire [7:0] soc_hdmi_out0_driver_sink_sink_payload_g;
wire [7:0] soc_hdmi_out0_driver_sink_sink_payload_b;
wire soc_hdmi_out0_driver_sink_sink_param_hsync;
wire soc_hdmi_out0_driver_sink_sink_param_vsync;
wire soc_hdmi_out0_driver_sink_sink_param_de;
wire hdmi_out0_pix_clk;
wire hdmi_out0_pix_rst;
wire hdmi_out0_pix5x_clk;
reg soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage_full = 1'd0;
wire soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage;
reg soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_re = 1'd0;
wire soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_read_re;
wire soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_read_r;
reg soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_read_w = 1'd0;
wire soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_write_re;
wire soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_write_r;
reg soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_write_w = 1'd0;
reg soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy_status = 1'd0;
reg [6:0] soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage_full = 7'd0;
wire [6:0] soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage;
reg soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_re = 1'd0;
reg [15:0] soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage_full = 16'd0;
wire [15:0] soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage;
reg soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_re = 1'd0;
wire [15:0] soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_r_status;
wire soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_locked;
wire soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_fb;
wire soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_clk0;
wire soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_clk1;
wire soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy;
wire [9:0] soc_hdmi_out0_driver_s7hdmioutclocking_data0;
wire [9:0] soc_hdmi_out0_driver_s7hdmioutclocking_data1;
reg soc_hdmi_out0_driver_s7hdmioutclocking_ce = 1'd0;
wire [1:0] soc_hdmi_out0_driver_s7hdmioutclocking_shift;
wire soc_hdmi_out0_driver_s7hdmioutclocking_pad_se;
reg [9:0] soc_hdmi_out0_driver_s7hdmioutclocking = 10'd31;
wire soc_hdmi_out0_driver_hdmi_phy_sink_valid;
wire soc_hdmi_out0_driver_hdmi_phy_sink_ready;
wire soc_hdmi_out0_driver_hdmi_phy_sink_first;
wire soc_hdmi_out0_driver_hdmi_phy_sink_last;
wire [7:0] soc_hdmi_out0_driver_hdmi_phy_sink_payload_r;
wire [7:0] soc_hdmi_out0_driver_hdmi_phy_sink_payload_g;
wire [7:0] soc_hdmi_out0_driver_hdmi_phy_sink_payload_b;
wire soc_hdmi_out0_driver_hdmi_phy_sink_param_hsync;
wire soc_hdmi_out0_driver_hdmi_phy_sink_param_vsync;
wire soc_hdmi_out0_driver_hdmi_phy_sink_param_de;
wire [7:0] soc_hdmi_out0_driver_hdmi_phy_es0_d0;
wire [1:0] soc_hdmi_out0_driver_hdmi_phy_es0_c;
wire soc_hdmi_out0_driver_hdmi_phy_es0_de;
reg [9:0] soc_hdmi_out0_driver_hdmi_phy_es0_out = 10'd0;
reg [7:0] soc_hdmi_out0_driver_hdmi_phy_es0_d1 = 8'd0;
reg [3:0] soc_hdmi_out0_driver_hdmi_phy_es0_n1d = 4'd0;
reg [8:0] soc_hdmi_out0_driver_hdmi_phy_es0_q_m = 9'd0;
wire soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n;
reg [8:0] soc_hdmi_out0_driver_hdmi_phy_es0_q_m_r = 9'd0;
reg [3:0] soc_hdmi_out0_driver_hdmi_phy_es0_n0q_m = 4'd0;
reg [3:0] soc_hdmi_out0_driver_hdmi_phy_es0_n1q_m = 4'd0;
reg signed [5:0] soc_hdmi_out0_driver_hdmi_phy_es0_cnt = 6'sd64;
reg [1:0] soc_hdmi_out0_driver_hdmi_phy_es0_new_c0 = 2'd0;
reg soc_hdmi_out0_driver_hdmi_phy_es0_new_de0 = 1'd0;
reg [1:0] soc_hdmi_out0_driver_hdmi_phy_es0_new_c1 = 2'd0;
reg soc_hdmi_out0_driver_hdmi_phy_es0_new_de1 = 1'd0;
reg [1:0] soc_hdmi_out0_driver_hdmi_phy_es0_new_c2 = 2'd0;
reg soc_hdmi_out0_driver_hdmi_phy_es0_new_de2 = 1'd0;
wire [9:0] soc_hdmi_out0_driver_hdmi_phy_es0_data;
reg soc_hdmi_out0_driver_hdmi_phy_es0_ce = 1'd0;
wire [1:0] soc_hdmi_out0_driver_hdmi_phy_es0_shift;
wire soc_hdmi_out0_driver_hdmi_phy_es0_pad_se;
wire [7:0] soc_hdmi_out0_driver_hdmi_phy_es1_d0;
wire [1:0] soc_hdmi_out0_driver_hdmi_phy_es1_c;
wire soc_hdmi_out0_driver_hdmi_phy_es1_de;
reg [9:0] soc_hdmi_out0_driver_hdmi_phy_es1_out = 10'd0;
reg [7:0] soc_hdmi_out0_driver_hdmi_phy_es1_d1 = 8'd0;
reg [3:0] soc_hdmi_out0_driver_hdmi_phy_es1_n1d = 4'd0;
reg [8:0] soc_hdmi_out0_driver_hdmi_phy_es1_q_m = 9'd0;
wire soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n;
reg [8:0] soc_hdmi_out0_driver_hdmi_phy_es1_q_m_r = 9'd0;
reg [3:0] soc_hdmi_out0_driver_hdmi_phy_es1_n0q_m = 4'd0;
reg [3:0] soc_hdmi_out0_driver_hdmi_phy_es1_n1q_m = 4'd0;
reg signed [5:0] soc_hdmi_out0_driver_hdmi_phy_es1_cnt = 6'sd64;
reg [1:0] soc_hdmi_out0_driver_hdmi_phy_es1_new_c0 = 2'd0;
reg soc_hdmi_out0_driver_hdmi_phy_es1_new_de0 = 1'd0;
reg [1:0] soc_hdmi_out0_driver_hdmi_phy_es1_new_c1 = 2'd0;
reg soc_hdmi_out0_driver_hdmi_phy_es1_new_de1 = 1'd0;
reg [1:0] soc_hdmi_out0_driver_hdmi_phy_es1_new_c2 = 2'd0;
reg soc_hdmi_out0_driver_hdmi_phy_es1_new_de2 = 1'd0;
wire [9:0] soc_hdmi_out0_driver_hdmi_phy_es1_data;
reg soc_hdmi_out0_driver_hdmi_phy_es1_ce = 1'd0;
wire [1:0] soc_hdmi_out0_driver_hdmi_phy_es1_shift;
wire soc_hdmi_out0_driver_hdmi_phy_es1_pad_se;
wire [7:0] soc_hdmi_out0_driver_hdmi_phy_es2_d0;
wire [1:0] soc_hdmi_out0_driver_hdmi_phy_es2_c;
wire soc_hdmi_out0_driver_hdmi_phy_es2_de;
reg [9:0] soc_hdmi_out0_driver_hdmi_phy_es2_out = 10'd0;
reg [7:0] soc_hdmi_out0_driver_hdmi_phy_es2_d1 = 8'd0;
reg [3:0] soc_hdmi_out0_driver_hdmi_phy_es2_n1d = 4'd0;
reg [8:0] soc_hdmi_out0_driver_hdmi_phy_es2_q_m = 9'd0;
wire soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n;
reg [8:0] soc_hdmi_out0_driver_hdmi_phy_es2_q_m_r = 9'd0;
reg [3:0] soc_hdmi_out0_driver_hdmi_phy_es2_n0q_m = 4'd0;
reg [3:0] soc_hdmi_out0_driver_hdmi_phy_es2_n1q_m = 4'd0;
reg signed [5:0] soc_hdmi_out0_driver_hdmi_phy_es2_cnt = 6'sd64;
reg [1:0] soc_hdmi_out0_driver_hdmi_phy_es2_new_c0 = 2'd0;
reg soc_hdmi_out0_driver_hdmi_phy_es2_new_de0 = 1'd0;
reg [1:0] soc_hdmi_out0_driver_hdmi_phy_es2_new_c1 = 2'd0;
reg soc_hdmi_out0_driver_hdmi_phy_es2_new_de1 = 1'd0;
reg [1:0] soc_hdmi_out0_driver_hdmi_phy_es2_new_c2 = 2'd0;
reg soc_hdmi_out0_driver_hdmi_phy_es2_new_de2 = 1'd0;
wire [9:0] soc_hdmi_out0_driver_hdmi_phy_es2_data;
reg soc_hdmi_out0_driver_hdmi_phy_es2_ce = 1'd0;
wire [1:0] soc_hdmi_out0_driver_hdmi_phy_es2_shift;
wire soc_hdmi_out0_driver_hdmi_phy_es2_pad_se;
wire soc_hdmi_out0_resetinserter_sink_sink_valid;
reg soc_hdmi_out0_resetinserter_sink_sink_ready = 1'd0;
wire [7:0] soc_hdmi_out0_resetinserter_sink_sink_payload_y;
wire [7:0] soc_hdmi_out0_resetinserter_sink_sink_payload_cb_cr;
wire soc_hdmi_out0_resetinserter_source_source_valid;
wire soc_hdmi_out0_resetinserter_source_source_ready;
reg soc_hdmi_out0_resetinserter_source_source_first = 1'd0;
reg soc_hdmi_out0_resetinserter_source_source_last = 1'd0;
wire [7:0] soc_hdmi_out0_resetinserter_source_source_payload_y;
wire [7:0] soc_hdmi_out0_resetinserter_source_source_payload_cb;
wire [7:0] soc_hdmi_out0_resetinserter_source_source_payload_cr;
reg soc_hdmi_out0_resetinserter_y_fifo_sink_valid = 1'd0;
wire soc_hdmi_out0_resetinserter_y_fifo_sink_ready;
reg soc_hdmi_out0_resetinserter_y_fifo_sink_first = 1'd0;
reg soc_hdmi_out0_resetinserter_y_fifo_sink_last = 1'd0;
reg [7:0] soc_hdmi_out0_resetinserter_y_fifo_sink_payload_data = 8'd0;
wire soc_hdmi_out0_resetinserter_y_fifo_source_valid;
wire soc_hdmi_out0_resetinserter_y_fifo_source_ready;
wire soc_hdmi_out0_resetinserter_y_fifo_source_first;
wire soc_hdmi_out0_resetinserter_y_fifo_source_last;
wire [7:0] soc_hdmi_out0_resetinserter_y_fifo_source_payload_data;
wire soc_hdmi_out0_resetinserter_y_fifo_syncfifo_we;
wire soc_hdmi_out0_resetinserter_y_fifo_syncfifo_writable;
wire soc_hdmi_out0_resetinserter_y_fifo_syncfifo_re;
wire soc_hdmi_out0_resetinserter_y_fifo_syncfifo_readable;
wire [9:0] soc_hdmi_out0_resetinserter_y_fifo_syncfifo_din;
wire [9:0] soc_hdmi_out0_resetinserter_y_fifo_syncfifo_dout;
reg [2:0] soc_hdmi_out0_resetinserter_y_fifo_level = 3'd0;
reg soc_hdmi_out0_resetinserter_y_fifo_replace = 1'd0;
reg [1:0] soc_hdmi_out0_resetinserter_y_fifo_produce = 2'd0;
reg [1:0] soc_hdmi_out0_resetinserter_y_fifo_consume = 2'd0;
reg [1:0] soc_hdmi_out0_resetinserter_y_fifo_wrport_adr = 2'd0;
wire [9:0] soc_hdmi_out0_resetinserter_y_fifo_wrport_dat_r;
wire soc_hdmi_out0_resetinserter_y_fifo_wrport_we;
wire [9:0] soc_hdmi_out0_resetinserter_y_fifo_wrport_dat_w;
wire soc_hdmi_out0_resetinserter_y_fifo_do_read;
wire [1:0] soc_hdmi_out0_resetinserter_y_fifo_rdport_adr;
wire [9:0] soc_hdmi_out0_resetinserter_y_fifo_rdport_dat_r;
wire [7:0] soc_hdmi_out0_resetinserter_y_fifo_fifo_in_payload_data;
wire soc_hdmi_out0_resetinserter_y_fifo_fifo_in_first;
wire soc_hdmi_out0_resetinserter_y_fifo_fifo_in_last;
wire [7:0] soc_hdmi_out0_resetinserter_y_fifo_fifo_out_payload_data;
wire soc_hdmi_out0_resetinserter_y_fifo_fifo_out_first;
wire soc_hdmi_out0_resetinserter_y_fifo_fifo_out_last;
reg soc_hdmi_out0_resetinserter_cb_fifo_sink_valid = 1'd0;
wire soc_hdmi_out0_resetinserter_cb_fifo_sink_ready;
reg soc_hdmi_out0_resetinserter_cb_fifo_sink_first = 1'd0;
reg soc_hdmi_out0_resetinserter_cb_fifo_sink_last = 1'd0;
reg [7:0] soc_hdmi_out0_resetinserter_cb_fifo_sink_payload_data = 8'd0;
wire soc_hdmi_out0_resetinserter_cb_fifo_source_valid;
wire soc_hdmi_out0_resetinserter_cb_fifo_source_ready;
wire soc_hdmi_out0_resetinserter_cb_fifo_source_first;
wire soc_hdmi_out0_resetinserter_cb_fifo_source_last;
wire [7:0] soc_hdmi_out0_resetinserter_cb_fifo_source_payload_data;
wire soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_we;
wire soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_writable;
wire soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_re;
wire soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_readable;
wire [9:0] soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_din;
wire [9:0] soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_dout;
reg [2:0] soc_hdmi_out0_resetinserter_cb_fifo_level = 3'd0;
reg soc_hdmi_out0_resetinserter_cb_fifo_replace = 1'd0;
reg [1:0] soc_hdmi_out0_resetinserter_cb_fifo_produce = 2'd0;
reg [1:0] soc_hdmi_out0_resetinserter_cb_fifo_consume = 2'd0;
reg [1:0] soc_hdmi_out0_resetinserter_cb_fifo_wrport_adr = 2'd0;
wire [9:0] soc_hdmi_out0_resetinserter_cb_fifo_wrport_dat_r;
wire soc_hdmi_out0_resetinserter_cb_fifo_wrport_we;
wire [9:0] soc_hdmi_out0_resetinserter_cb_fifo_wrport_dat_w;
wire soc_hdmi_out0_resetinserter_cb_fifo_do_read;
wire [1:0] soc_hdmi_out0_resetinserter_cb_fifo_rdport_adr;
wire [9:0] soc_hdmi_out0_resetinserter_cb_fifo_rdport_dat_r;
wire [7:0] soc_hdmi_out0_resetinserter_cb_fifo_fifo_in_payload_data;
wire soc_hdmi_out0_resetinserter_cb_fifo_fifo_in_first;
wire soc_hdmi_out0_resetinserter_cb_fifo_fifo_in_last;
wire [7:0] soc_hdmi_out0_resetinserter_cb_fifo_fifo_out_payload_data;
wire soc_hdmi_out0_resetinserter_cb_fifo_fifo_out_first;
wire soc_hdmi_out0_resetinserter_cb_fifo_fifo_out_last;
reg soc_hdmi_out0_resetinserter_cr_fifo_sink_valid = 1'd0;
wire soc_hdmi_out0_resetinserter_cr_fifo_sink_ready;
reg soc_hdmi_out0_resetinserter_cr_fifo_sink_first = 1'd0;
reg soc_hdmi_out0_resetinserter_cr_fifo_sink_last = 1'd0;
reg [7:0] soc_hdmi_out0_resetinserter_cr_fifo_sink_payload_data = 8'd0;
wire soc_hdmi_out0_resetinserter_cr_fifo_source_valid;
wire soc_hdmi_out0_resetinserter_cr_fifo_source_ready;
wire soc_hdmi_out0_resetinserter_cr_fifo_source_first;
wire soc_hdmi_out0_resetinserter_cr_fifo_source_last;
wire [7:0] soc_hdmi_out0_resetinserter_cr_fifo_source_payload_data;
wire soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_we;
wire soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_writable;
wire soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_re;
wire soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_readable;
wire [9:0] soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_din;
wire [9:0] soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_dout;
reg [2:0] soc_hdmi_out0_resetinserter_cr_fifo_level = 3'd0;
reg soc_hdmi_out0_resetinserter_cr_fifo_replace = 1'd0;
reg [1:0] soc_hdmi_out0_resetinserter_cr_fifo_produce = 2'd0;
reg [1:0] soc_hdmi_out0_resetinserter_cr_fifo_consume = 2'd0;
reg [1:0] soc_hdmi_out0_resetinserter_cr_fifo_wrport_adr = 2'd0;
wire [9:0] soc_hdmi_out0_resetinserter_cr_fifo_wrport_dat_r;
wire soc_hdmi_out0_resetinserter_cr_fifo_wrport_we;
wire [9:0] soc_hdmi_out0_resetinserter_cr_fifo_wrport_dat_w;
wire soc_hdmi_out0_resetinserter_cr_fifo_do_read;
wire [1:0] soc_hdmi_out0_resetinserter_cr_fifo_rdport_adr;
wire [9:0] soc_hdmi_out0_resetinserter_cr_fifo_rdport_dat_r;
wire [7:0] soc_hdmi_out0_resetinserter_cr_fifo_fifo_in_payload_data;
wire soc_hdmi_out0_resetinserter_cr_fifo_fifo_in_first;
wire soc_hdmi_out0_resetinserter_cr_fifo_fifo_in_last;
wire [7:0] soc_hdmi_out0_resetinserter_cr_fifo_fifo_out_payload_data;
wire soc_hdmi_out0_resetinserter_cr_fifo_fifo_out_first;
wire soc_hdmi_out0_resetinserter_cr_fifo_fifo_out_last;
reg soc_hdmi_out0_resetinserter_parity_in = 1'd0;
reg soc_hdmi_out0_resetinserter_parity_out = 1'd0;
wire soc_hdmi_out0_resetinserter_reset;
wire soc_hdmi_out0_sink_valid;
wire soc_hdmi_out0_sink_ready;
wire soc_hdmi_out0_sink_first;
wire soc_hdmi_out0_sink_last;
wire [7:0] soc_hdmi_out0_sink_payload_y;
wire [7:0] soc_hdmi_out0_sink_payload_cb;
wire [7:0] soc_hdmi_out0_sink_payload_cr;
wire soc_hdmi_out0_source_valid;
wire soc_hdmi_out0_source_ready;
wire soc_hdmi_out0_source_first;
wire soc_hdmi_out0_source_last;
wire [7:0] soc_hdmi_out0_source_payload_r;
wire [7:0] soc_hdmi_out0_source_payload_g;
wire [7:0] soc_hdmi_out0_source_payload_b;
wire [7:0] soc_hdmi_out0_sink_y;
wire [7:0] soc_hdmi_out0_sink_cb;
wire [7:0] soc_hdmi_out0_sink_cr;
reg [7:0] soc_hdmi_out0_source_r = 8'd0;
reg [7:0] soc_hdmi_out0_source_g = 8'd0;
reg [7:0] soc_hdmi_out0_source_b = 8'd0;
reg [7:0] soc_hdmi_out0_record0_ycbcr_n_y = 8'd0;
reg [7:0] soc_hdmi_out0_record0_ycbcr_n_cb = 8'd0;
reg [7:0] soc_hdmi_out0_record0_ycbcr_n_cr = 8'd0;
reg [7:0] soc_hdmi_out0_record1_ycbcr_n_y = 8'd0;
reg [7:0] soc_hdmi_out0_record1_ycbcr_n_cb = 8'd0;
reg [7:0] soc_hdmi_out0_record1_ycbcr_n_cr = 8'd0;
reg [7:0] soc_hdmi_out0_record2_ycbcr_n_y = 8'd0;
reg [7:0] soc_hdmi_out0_record2_ycbcr_n_cb = 8'd0;
reg [7:0] soc_hdmi_out0_record2_ycbcr_n_cr = 8'd0;
reg [7:0] soc_hdmi_out0_record3_ycbcr_n_y = 8'd0;
reg [7:0] soc_hdmi_out0_record3_ycbcr_n_cb = 8'd0;
reg [7:0] soc_hdmi_out0_record3_ycbcr_n_cr = 8'd0;
reg signed [8:0] soc_hdmi_out0_cb_minus_coffset = 9'sd512;
reg signed [8:0] soc_hdmi_out0_cr_minus_coffset = 9'sd512;
reg signed [8:0] soc_hdmi_out0_y_minus_yoffset = 9'sd512;
reg signed [19:0] soc_hdmi_out0_cr_minus_coffset_mult_acoef = 20'sd1048576;
reg signed [19:0] soc_hdmi_out0_cb_minus_coffset_mult_bcoef = 20'sd1048576;
reg signed [19:0] soc_hdmi_out0_cr_minus_coffset_mult_ccoef = 20'sd1048576;
reg signed [19:0] soc_hdmi_out0_cb_minus_coffset_mult_dcoef = 20'sd1048576;
reg signed [11:0] soc_hdmi_out0_r = 12'sd4096;
reg signed [11:0] soc_hdmi_out0_g = 12'sd4096;
reg signed [11:0] soc_hdmi_out0_b = 12'sd4096;
wire soc_hdmi_out0_ce;
wire soc_hdmi_out0_pipe_ce;
wire soc_hdmi_out0_busy;
reg soc_hdmi_out0_valid_n0 = 1'd0;
reg soc_hdmi_out0_valid_n1 = 1'd0;
reg soc_hdmi_out0_valid_n2 = 1'd0;
reg soc_hdmi_out0_valid_n3 = 1'd0;
reg soc_hdmi_out0_first_n0 = 1'd0;
reg soc_hdmi_out0_last_n0 = 1'd0;
reg soc_hdmi_out0_first_n1 = 1'd0;
reg soc_hdmi_out0_last_n1 = 1'd0;
reg soc_hdmi_out0_first_n2 = 1'd0;
reg soc_hdmi_out0_last_n2 = 1'd0;
reg soc_hdmi_out0_first_n3 = 1'd0;
reg soc_hdmi_out0_last_n3 = 1'd0;
wire soc_hdmi_out0_sink_payload_hsync;
wire soc_hdmi_out0_sink_payload_vsync;
wire soc_hdmi_out0_sink_payload_de;
wire soc_hdmi_out0_source_payload_hsync;
wire soc_hdmi_out0_source_payload_vsync;
wire soc_hdmi_out0_source_payload_de;
reg soc_hdmi_out0_next_s0 = 1'd0;
reg soc_hdmi_out0_next_s1 = 1'd0;
reg soc_hdmi_out0_next_s2 = 1'd0;
reg soc_hdmi_out0_next_s3 = 1'd0;
reg soc_hdmi_out0_next_s4 = 1'd0;
reg soc_hdmi_out0_next_s5 = 1'd0;
reg soc_hdmi_out0_next_s6 = 1'd0;
reg soc_hdmi_out0_next_s7 = 1'd0;
reg soc_hdmi_out0_next_s8 = 1'd0;
reg soc_hdmi_out0_next_s9 = 1'd0;
reg soc_hdmi_out0_next_s10 = 1'd0;
reg soc_hdmi_out0_next_s11 = 1'd0;
reg soc_hdmi_out0_next_s12 = 1'd0;
reg soc_hdmi_out0_next_s13 = 1'd0;
reg soc_hdmi_out0_next_s14 = 1'd0;
reg soc_hdmi_out0_next_s15 = 1'd0;
reg soc_hdmi_out0_next_s16 = 1'd0;
reg soc_hdmi_out0_next_s17 = 1'd0;
reg soc_hdmi_out0_de_r = 1'd0;
reg soc_hdmi_out0_core_source_valid_d = 1'd0;
reg [15:0] soc_hdmi_out0_core_source_data_d = 16'd0;
reg [2:0] vns_wishbonestreamingbridge_state = 3'd0;
reg [2:0] vns_wishbonestreamingbridge_next_state = 3'd0;
reg [1:0] vns_oled_state = 2'd0;
reg [1:0] vns_oled_next_state = 2'd0;
reg [1:0] vns_refresher_state = 2'd0;
reg [1:0] vns_refresher_next_state = 2'd0;
reg [2:0] vns_bankmachine0_state = 3'd0;
reg [2:0] vns_bankmachine0_next_state = 3'd0;
reg [2:0] vns_bankmachine1_state = 3'd0;
reg [2:0] vns_bankmachine1_next_state = 3'd0;
reg [2:0] vns_bankmachine2_state = 3'd0;
reg [2:0] vns_bankmachine2_next_state = 3'd0;
reg [2:0] vns_bankmachine3_state = 3'd0;
reg [2:0] vns_bankmachine3_next_state = 3'd0;
reg [2:0] vns_bankmachine4_state = 3'd0;
reg [2:0] vns_bankmachine4_next_state = 3'd0;
reg [2:0] vns_bankmachine5_state = 3'd0;
reg [2:0] vns_bankmachine5_next_state = 3'd0;
reg [2:0] vns_bankmachine6_state = 3'd0;
reg [2:0] vns_bankmachine6_next_state = 3'd0;
reg [2:0] vns_bankmachine7_state = 3'd0;
reg [2:0] vns_bankmachine7_next_state = 3'd0;
reg [3:0] vns_multiplexer_state = 4'd0;
reg [3:0] vns_multiplexer_next_state = 4'd0;
wire [2:0] vns_cba0;
wire [21:0] vns_rca0;
wire [2:0] vns_cba1;
wire [21:0] vns_rca1;
wire [2:0] vns_cba2;
wire [21:0] vns_rca2;
wire [2:0] vns_roundrobin0_request;
reg [1:0] vns_roundrobin0_grant = 2'd0;
wire vns_roundrobin0_ce;
wire [2:0] vns_roundrobin1_request;
reg [1:0] vns_roundrobin1_grant = 2'd0;
wire vns_roundrobin1_ce;
wire [2:0] vns_roundrobin2_request;
reg [1:0] vns_roundrobin2_grant = 2'd0;
wire vns_roundrobin2_ce;
wire [2:0] vns_roundrobin3_request;
reg [1:0] vns_roundrobin3_grant = 2'd0;
wire vns_roundrobin3_ce;
wire [2:0] vns_roundrobin4_request;
reg [1:0] vns_roundrobin4_grant = 2'd0;
wire vns_roundrobin4_ce;
wire [2:0] vns_roundrobin5_request;
reg [1:0] vns_roundrobin5_grant = 2'd0;
wire vns_roundrobin5_ce;
wire [2:0] vns_roundrobin6_request;
reg [1:0] vns_roundrobin6_grant = 2'd0;
wire vns_roundrobin6_ce;
wire [2:0] vns_roundrobin7_request;
reg [1:0] vns_roundrobin7_grant = 2'd0;
wire vns_roundrobin7_ce;
reg vns_new_master_wdata_ready0 = 1'd0;
reg vns_new_master_wdata_ready1 = 1'd0;
reg vns_new_master_wdata_ready2 = 1'd0;
reg vns_new_master_wdata_ready3 = 1'd0;
reg vns_new_master_wdata_ready4 = 1'd0;
reg vns_new_master_wdata_ready5 = 1'd0;
reg vns_new_master_wdata_ready6 = 1'd0;
reg vns_new_master_wdata_ready7 = 1'd0;
reg vns_new_master_wdata_ready8 = 1'd0;
reg vns_new_master_rdata_valid0 = 1'd0;
reg vns_new_master_rdata_valid1 = 1'd0;
reg vns_new_master_rdata_valid2 = 1'd0;
reg vns_new_master_rdata_valid3 = 1'd0;
reg vns_new_master_rdata_valid4 = 1'd0;
reg vns_new_master_rdata_valid5 = 1'd0;
reg vns_new_master_rdata_valid6 = 1'd0;
reg vns_new_master_rdata_valid7 = 1'd0;
reg vns_new_master_rdata_valid8 = 1'd0;
reg vns_new_master_rdata_valid9 = 1'd0;
reg vns_new_master_rdata_valid10 = 1'd0;
reg vns_new_master_rdata_valid11 = 1'd0;
reg vns_new_master_rdata_valid12 = 1'd0;
reg vns_new_master_rdata_valid13 = 1'd0;
reg vns_new_master_rdata_valid14 = 1'd0;
reg vns_new_master_rdata_valid15 = 1'd0;
reg vns_new_master_rdata_valid16 = 1'd0;
reg vns_new_master_rdata_valid17 = 1'd0;
reg vns_new_master_rdata_valid18 = 1'd0;
reg vns_new_master_rdata_valid19 = 1'd0;
reg vns_new_master_rdata_valid20 = 1'd0;
reg [2:0] vns_fullmemorywe_state = 3'd0;
reg [2:0] vns_fullmemorywe_next_state = 3'd0;
reg [1:0] vns_litedramwishbonebridge_state = 2'd0;
reg [1:0] vns_litedramwishbonebridge_next_state = 2'd0;
reg vns_clockdomainsrenamer0_state = 1'd0;
reg vns_clockdomainsrenamer0_next_state = 1'd0;
reg vns_clockdomainsrenamer1_state = 1'd0;
reg vns_clockdomainsrenamer1_next_state = 1'd0;
reg [1:0] vns_clockdomainsrenamer2_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer2_next_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer3_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer3_next_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer4_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer4_next_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer5_state = 2'd0;
reg [1:0] vns_clockdomainsrenamer5_next_state = 2'd0;
reg vns_clockdomainsrenamer6_state = 1'd0;
reg vns_clockdomainsrenamer6_next_state = 1'd0;
reg [1:0] vns_liteethmacsramwriter_state = 2'd0;
reg [1:0] vns_liteethmacsramwriter_next_state = 2'd0;
reg [1:0] vns_liteethmacsramreader_state = 2'd0;
reg [1:0] vns_liteethmacsramreader_next_state = 2'd0;
reg [3:0] vns_edid_state = 4'd0;
reg [3:0] vns_edid_next_state = 4'd0;
reg [1:0] vns_dma_state = 2'd0;
reg [1:0] vns_dma_next_state = 2'd0;
reg vns_videoout_state = 1'd0;
reg vns_videoout_next_state = 1'd0;
reg [27:0] soc_hdmi_out0_core_dmareader_offset_next_value = 28'd0;
reg soc_hdmi_out0_core_dmareader_offset_next_value_ce = 1'd0;
wire vns_wb_sdram_con_request;
wire vns_wb_sdram_con_grant;
wire [29:0] vns_videosoc_shared_adr;
wire [31:0] vns_videosoc_shared_dat_w;
wire [31:0] vns_videosoc_shared_dat_r;
wire [3:0] vns_videosoc_shared_sel;
wire vns_videosoc_shared_cyc;
wire vns_videosoc_shared_stb;
wire vns_videosoc_shared_ack;
wire vns_videosoc_shared_we;
wire [2:0] vns_videosoc_shared_cti;
wire [1:0] vns_videosoc_shared_bte;
wire vns_videosoc_shared_err;
wire [2:0] vns_videosoc_request;
reg [1:0] vns_videosoc_grant = 2'd0;
reg [5:0] vns_videosoc_slave_sel = 6'd0;
reg [5:0] vns_videosoc_slave_sel_r = 6'd0;
wire [13:0] vns_videosoc_interface0_bank_bus_adr;
wire vns_videosoc_interface0_bank_bus_we;
wire [7:0] vns_videosoc_interface0_bank_bus_dat_w;
reg [7:0] vns_videosoc_interface0_bank_bus_dat_r = 8'd0;
wire vns_videosoc_csrbank0_dly_sel0_re;
wire [1:0] vns_videosoc_csrbank0_dly_sel0_r;
wire [1:0] vns_videosoc_csrbank0_dly_sel0_w;
wire vns_videosoc_csrbank0_sel;
wire [13:0] vns_videosoc_interface1_bank_bus_adr;
wire vns_videosoc_interface1_bank_bus_we;
wire [7:0] vns_videosoc_interface1_bank_bus_dat_w;
reg [7:0] vns_videosoc_interface1_bank_bus_dat_r = 8'd0;
wire vns_videosoc_csrbank1_sram_writer_slot_re;
wire vns_videosoc_csrbank1_sram_writer_slot_r;
wire vns_videosoc_csrbank1_sram_writer_slot_w;
wire vns_videosoc_csrbank1_sram_writer_length3_re;
wire [7:0] vns_videosoc_csrbank1_sram_writer_length3_r;
wire [7:0] vns_videosoc_csrbank1_sram_writer_length3_w;
wire vns_videosoc_csrbank1_sram_writer_length2_re;
wire [7:0] vns_videosoc_csrbank1_sram_writer_length2_r;
wire [7:0] vns_videosoc_csrbank1_sram_writer_length2_w;
wire vns_videosoc_csrbank1_sram_writer_length1_re;
wire [7:0] vns_videosoc_csrbank1_sram_writer_length1_r;
wire [7:0] vns_videosoc_csrbank1_sram_writer_length1_w;
wire vns_videosoc_csrbank1_sram_writer_length0_re;
wire [7:0] vns_videosoc_csrbank1_sram_writer_length0_r;
wire [7:0] vns_videosoc_csrbank1_sram_writer_length0_w;
wire vns_videosoc_csrbank1_sram_writer_ev_enable0_re;
wire vns_videosoc_csrbank1_sram_writer_ev_enable0_r;
wire vns_videosoc_csrbank1_sram_writer_ev_enable0_w;
wire vns_videosoc_csrbank1_sram_reader_ready_re;
wire vns_videosoc_csrbank1_sram_reader_ready_r;
wire vns_videosoc_csrbank1_sram_reader_ready_w;
wire vns_videosoc_csrbank1_sram_reader_slot0_re;
wire vns_videosoc_csrbank1_sram_reader_slot0_r;
wire vns_videosoc_csrbank1_sram_reader_slot0_w;
wire vns_videosoc_csrbank1_sram_reader_length1_re;
wire [2:0] vns_videosoc_csrbank1_sram_reader_length1_r;
wire [2:0] vns_videosoc_csrbank1_sram_reader_length1_w;
wire vns_videosoc_csrbank1_sram_reader_length0_re;
wire [7:0] vns_videosoc_csrbank1_sram_reader_length0_r;
wire [7:0] vns_videosoc_csrbank1_sram_reader_length0_w;
wire vns_videosoc_csrbank1_sram_reader_ev_enable0_re;
wire vns_videosoc_csrbank1_sram_reader_ev_enable0_r;
wire vns_videosoc_csrbank1_sram_reader_ev_enable0_w;
wire vns_videosoc_csrbank1_preamble_crc_re;
wire vns_videosoc_csrbank1_preamble_crc_r;
wire vns_videosoc_csrbank1_preamble_crc_w;
wire vns_videosoc_csrbank1_sel;
wire [13:0] vns_videosoc_interface2_bank_bus_adr;
wire vns_videosoc_interface2_bank_bus_we;
wire [7:0] vns_videosoc_interface2_bank_bus_dat_w;
reg [7:0] vns_videosoc_interface2_bank_bus_dat_r = 8'd0;
wire vns_videosoc_csrbank2_crg_reset0_re;
wire vns_videosoc_csrbank2_crg_reset0_r;
wire vns_videosoc_csrbank2_crg_reset0_w;
wire vns_videosoc_csrbank2_mdio_w0_re;
wire [2:0] vns_videosoc_csrbank2_mdio_w0_r;
wire [2:0] vns_videosoc_csrbank2_mdio_w0_w;
wire vns_videosoc_csrbank2_mdio_r_re;
wire vns_videosoc_csrbank2_mdio_r_r;
wire vns_videosoc_csrbank2_mdio_r_w;
wire vns_videosoc_csrbank2_sel;
wire [13:0] vns_videosoc_sram_bus_adr;
wire vns_videosoc_sram_bus_we;
wire [7:0] vns_videosoc_sram_bus_dat_w;
reg [7:0] vns_videosoc_sram_bus_dat_r = 8'd0;
wire [6:0] vns_videosoc_adr;
wire [7:0] vns_videosoc_dat_r;
wire vns_videosoc_we;
wire [7:0] vns_videosoc_dat_w;
wire vns_videosoc_sel;
reg vns_videosoc_sel_r = 1'd0;
wire [13:0] vns_videosoc_interface3_bank_bus_adr;
wire vns_videosoc_interface3_bank_bus_we;
wire [7:0] vns_videosoc_interface3_bank_bus_dat_w;
reg [7:0] vns_videosoc_interface3_bank_bus_dat_r = 8'd0;
wire vns_videosoc_csrbank3_edid_hpd_notif_re;
wire vns_videosoc_csrbank3_edid_hpd_notif_r;
wire vns_videosoc_csrbank3_edid_hpd_notif_w;
wire vns_videosoc_csrbank3_edid_hpd_en0_re;
wire vns_videosoc_csrbank3_edid_hpd_en0_r;
wire vns_videosoc_csrbank3_edid_hpd_en0_w;
wire vns_videosoc_csrbank3_clocking_mmcm_reset0_re;
wire vns_videosoc_csrbank3_clocking_mmcm_reset0_r;
wire vns_videosoc_csrbank3_clocking_mmcm_reset0_w;
wire vns_videosoc_csrbank3_clocking_locked_re;
wire vns_videosoc_csrbank3_clocking_locked_r;
wire vns_videosoc_csrbank3_clocking_locked_w;
wire vns_videosoc_csrbank3_clocking_mmcm_drdy_re;
wire vns_videosoc_csrbank3_clocking_mmcm_drdy_r;
wire vns_videosoc_csrbank3_clocking_mmcm_drdy_w;
wire vns_videosoc_csrbank3_clocking_mmcm_adr0_re;
wire [6:0] vns_videosoc_csrbank3_clocking_mmcm_adr0_r;
wire [6:0] vns_videosoc_csrbank3_clocking_mmcm_adr0_w;
wire vns_videosoc_csrbank3_clocking_mmcm_dat_w1_re;
wire [7:0] vns_videosoc_csrbank3_clocking_mmcm_dat_w1_r;
wire [7:0] vns_videosoc_csrbank3_clocking_mmcm_dat_w1_w;
wire vns_videosoc_csrbank3_clocking_mmcm_dat_w0_re;
wire [7:0] vns_videosoc_csrbank3_clocking_mmcm_dat_w0_r;
wire [7:0] vns_videosoc_csrbank3_clocking_mmcm_dat_w0_w;
wire vns_videosoc_csrbank3_clocking_mmcm_dat_r1_re;
wire [7:0] vns_videosoc_csrbank3_clocking_mmcm_dat_r1_r;
wire [7:0] vns_videosoc_csrbank3_clocking_mmcm_dat_r1_w;
wire vns_videosoc_csrbank3_clocking_mmcm_dat_r0_re;
wire [7:0] vns_videosoc_csrbank3_clocking_mmcm_dat_r0_r;
wire [7:0] vns_videosoc_csrbank3_clocking_mmcm_dat_r0_w;
wire vns_videosoc_csrbank3_data0_cap_phase_re;
wire [1:0] vns_videosoc_csrbank3_data0_cap_phase_r;
wire [1:0] vns_videosoc_csrbank3_data0_cap_phase_w;
wire vns_videosoc_csrbank3_data0_charsync_char_synced_re;
wire vns_videosoc_csrbank3_data0_charsync_char_synced_r;
wire vns_videosoc_csrbank3_data0_charsync_char_synced_w;
wire vns_videosoc_csrbank3_data0_charsync_ctl_pos_re;
wire [3:0] vns_videosoc_csrbank3_data0_charsync_ctl_pos_r;
wire [3:0] vns_videosoc_csrbank3_data0_charsync_ctl_pos_w;
wire vns_videosoc_csrbank3_data0_wer_value2_re;
wire [7:0] vns_videosoc_csrbank3_data0_wer_value2_r;
wire [7:0] vns_videosoc_csrbank3_data0_wer_value2_w;
wire vns_videosoc_csrbank3_data0_wer_value1_re;
wire [7:0] vns_videosoc_csrbank3_data0_wer_value1_r;
wire [7:0] vns_videosoc_csrbank3_data0_wer_value1_w;
wire vns_videosoc_csrbank3_data0_wer_value0_re;
wire [7:0] vns_videosoc_csrbank3_data0_wer_value0_r;
wire [7:0] vns_videosoc_csrbank3_data0_wer_value0_w;
wire vns_videosoc_csrbank3_data1_cap_phase_re;
wire [1:0] vns_videosoc_csrbank3_data1_cap_phase_r;
wire [1:0] vns_videosoc_csrbank3_data1_cap_phase_w;
wire vns_videosoc_csrbank3_data1_charsync_char_synced_re;
wire vns_videosoc_csrbank3_data1_charsync_char_synced_r;
wire vns_videosoc_csrbank3_data1_charsync_char_synced_w;
wire vns_videosoc_csrbank3_data1_charsync_ctl_pos_re;
wire [3:0] vns_videosoc_csrbank3_data1_charsync_ctl_pos_r;
wire [3:0] vns_videosoc_csrbank3_data1_charsync_ctl_pos_w;
wire vns_videosoc_csrbank3_data1_wer_value2_re;
wire [7:0] vns_videosoc_csrbank3_data1_wer_value2_r;
wire [7:0] vns_videosoc_csrbank3_data1_wer_value2_w;
wire vns_videosoc_csrbank3_data1_wer_value1_re;
wire [7:0] vns_videosoc_csrbank3_data1_wer_value1_r;
wire [7:0] vns_videosoc_csrbank3_data1_wer_value1_w;
wire vns_videosoc_csrbank3_data1_wer_value0_re;
wire [7:0] vns_videosoc_csrbank3_data1_wer_value0_r;
wire [7:0] vns_videosoc_csrbank3_data1_wer_value0_w;
wire vns_videosoc_csrbank3_data2_cap_phase_re;
wire [1:0] vns_videosoc_csrbank3_data2_cap_phase_r;
wire [1:0] vns_videosoc_csrbank3_data2_cap_phase_w;
wire vns_videosoc_csrbank3_data2_charsync_char_synced_re;
wire vns_videosoc_csrbank3_data2_charsync_char_synced_r;
wire vns_videosoc_csrbank3_data2_charsync_char_synced_w;
wire vns_videosoc_csrbank3_data2_charsync_ctl_pos_re;
wire [3:0] vns_videosoc_csrbank3_data2_charsync_ctl_pos_r;
wire [3:0] vns_videosoc_csrbank3_data2_charsync_ctl_pos_w;
wire vns_videosoc_csrbank3_data2_wer_value2_re;
wire [7:0] vns_videosoc_csrbank3_data2_wer_value2_r;
wire [7:0] vns_videosoc_csrbank3_data2_wer_value2_w;
wire vns_videosoc_csrbank3_data2_wer_value1_re;
wire [7:0] vns_videosoc_csrbank3_data2_wer_value1_r;
wire [7:0] vns_videosoc_csrbank3_data2_wer_value1_w;
wire vns_videosoc_csrbank3_data2_wer_value0_re;
wire [7:0] vns_videosoc_csrbank3_data2_wer_value0_r;
wire [7:0] vns_videosoc_csrbank3_data2_wer_value0_w;
wire vns_videosoc_csrbank3_chansync_channels_synced_re;
wire vns_videosoc_csrbank3_chansync_channels_synced_r;
wire vns_videosoc_csrbank3_chansync_channels_synced_w;
wire vns_videosoc_csrbank3_resdetection_hres1_re;
wire [2:0] vns_videosoc_csrbank3_resdetection_hres1_r;
wire [2:0] vns_videosoc_csrbank3_resdetection_hres1_w;
wire vns_videosoc_csrbank3_resdetection_hres0_re;
wire [7:0] vns_videosoc_csrbank3_resdetection_hres0_r;
wire [7:0] vns_videosoc_csrbank3_resdetection_hres0_w;
wire vns_videosoc_csrbank3_resdetection_vres1_re;
wire [2:0] vns_videosoc_csrbank3_resdetection_vres1_r;
wire [2:0] vns_videosoc_csrbank3_resdetection_vres1_w;
wire vns_videosoc_csrbank3_resdetection_vres0_re;
wire [7:0] vns_videosoc_csrbank3_resdetection_vres0_r;
wire [7:0] vns_videosoc_csrbank3_resdetection_vres0_w;
wire vns_videosoc_csrbank3_dma_frame_size3_re;
wire [4:0] vns_videosoc_csrbank3_dma_frame_size3_r;
wire [4:0] vns_videosoc_csrbank3_dma_frame_size3_w;
wire vns_videosoc_csrbank3_dma_frame_size2_re;
wire [7:0] vns_videosoc_csrbank3_dma_frame_size2_r;
wire [7:0] vns_videosoc_csrbank3_dma_frame_size2_w;
wire vns_videosoc_csrbank3_dma_frame_size1_re;
wire [7:0] vns_videosoc_csrbank3_dma_frame_size1_r;
wire [7:0] vns_videosoc_csrbank3_dma_frame_size1_w;
wire vns_videosoc_csrbank3_dma_frame_size0_re;
wire [7:0] vns_videosoc_csrbank3_dma_frame_size0_r;
wire [7:0] vns_videosoc_csrbank3_dma_frame_size0_w;
wire vns_videosoc_csrbank3_dma_slot0_status0_re;
wire [1:0] vns_videosoc_csrbank3_dma_slot0_status0_r;
wire [1:0] vns_videosoc_csrbank3_dma_slot0_status0_w;
wire vns_videosoc_csrbank3_dma_slot0_address3_re;
wire [4:0] vns_videosoc_csrbank3_dma_slot0_address3_r;
wire [4:0] vns_videosoc_csrbank3_dma_slot0_address3_w;
wire vns_videosoc_csrbank3_dma_slot0_address2_re;
wire [7:0] vns_videosoc_csrbank3_dma_slot0_address2_r;
wire [7:0] vns_videosoc_csrbank3_dma_slot0_address2_w;
wire vns_videosoc_csrbank3_dma_slot0_address1_re;
wire [7:0] vns_videosoc_csrbank3_dma_slot0_address1_r;
wire [7:0] vns_videosoc_csrbank3_dma_slot0_address1_w;
wire vns_videosoc_csrbank3_dma_slot0_address0_re;
wire [7:0] vns_videosoc_csrbank3_dma_slot0_address0_r;
wire [7:0] vns_videosoc_csrbank3_dma_slot0_address0_w;
wire vns_videosoc_csrbank3_dma_slot1_status0_re;
wire [1:0] vns_videosoc_csrbank3_dma_slot1_status0_r;
wire [1:0] vns_videosoc_csrbank3_dma_slot1_status0_w;
wire vns_videosoc_csrbank3_dma_slot1_address3_re;
wire [4:0] vns_videosoc_csrbank3_dma_slot1_address3_r;
wire [4:0] vns_videosoc_csrbank3_dma_slot1_address3_w;
wire vns_videosoc_csrbank3_dma_slot1_address2_re;
wire [7:0] vns_videosoc_csrbank3_dma_slot1_address2_r;
wire [7:0] vns_videosoc_csrbank3_dma_slot1_address2_w;
wire vns_videosoc_csrbank3_dma_slot1_address1_re;
wire [7:0] vns_videosoc_csrbank3_dma_slot1_address1_r;
wire [7:0] vns_videosoc_csrbank3_dma_slot1_address1_w;
wire vns_videosoc_csrbank3_dma_slot1_address0_re;
wire [7:0] vns_videosoc_csrbank3_dma_slot1_address0_r;
wire [7:0] vns_videosoc_csrbank3_dma_slot1_address0_w;
wire vns_videosoc_csrbank3_dma_ev_enable0_re;
wire [1:0] vns_videosoc_csrbank3_dma_ev_enable0_r;
wire [1:0] vns_videosoc_csrbank3_dma_ev_enable0_w;
wire vns_videosoc_csrbank3_sel;
wire [13:0] vns_videosoc_interface4_bank_bus_adr;
wire vns_videosoc_interface4_bank_bus_we;
wire [7:0] vns_videosoc_interface4_bank_bus_dat_w;
reg [7:0] vns_videosoc_interface4_bank_bus_dat_r = 8'd0;
wire vns_videosoc_csrbank4_value3_re;
wire [7:0] vns_videosoc_csrbank4_value3_r;
wire [7:0] vns_videosoc_csrbank4_value3_w;
wire vns_videosoc_csrbank4_value2_re;
wire [7:0] vns_videosoc_csrbank4_value2_r;
wire [7:0] vns_videosoc_csrbank4_value2_w;
wire vns_videosoc_csrbank4_value1_re;
wire [7:0] vns_videosoc_csrbank4_value1_r;
wire [7:0] vns_videosoc_csrbank4_value1_w;
wire vns_videosoc_csrbank4_value0_re;
wire [7:0] vns_videosoc_csrbank4_value0_r;
wire [7:0] vns_videosoc_csrbank4_value0_w;
wire vns_videosoc_csrbank4_sel;
wire [13:0] vns_videosoc_interface5_bank_bus_adr;
wire vns_videosoc_interface5_bank_bus_we;
wire [7:0] vns_videosoc_interface5_bank_bus_dat_w;
reg [7:0] vns_videosoc_interface5_bank_bus_dat_r = 8'd0;
wire vns_videosoc_csrbank5_core_underflow_enable0_re;
wire vns_videosoc_csrbank5_core_underflow_enable0_r;
wire vns_videosoc_csrbank5_core_underflow_enable0_w;
wire vns_videosoc_csrbank5_core_underflow_counter3_re;
wire [7:0] vns_videosoc_csrbank5_core_underflow_counter3_r;
wire [7:0] vns_videosoc_csrbank5_core_underflow_counter3_w;
wire vns_videosoc_csrbank5_core_underflow_counter2_re;
wire [7:0] vns_videosoc_csrbank5_core_underflow_counter2_r;
wire [7:0] vns_videosoc_csrbank5_core_underflow_counter2_w;
wire vns_videosoc_csrbank5_core_underflow_counter1_re;
wire [7:0] vns_videosoc_csrbank5_core_underflow_counter1_r;
wire [7:0] vns_videosoc_csrbank5_core_underflow_counter1_w;
wire vns_videosoc_csrbank5_core_underflow_counter0_re;
wire [7:0] vns_videosoc_csrbank5_core_underflow_counter0_r;
wire [7:0] vns_videosoc_csrbank5_core_underflow_counter0_w;
wire vns_videosoc_csrbank5_core_initiator_enable0_re;
wire vns_videosoc_csrbank5_core_initiator_enable0_r;
wire vns_videosoc_csrbank5_core_initiator_enable0_w;
reg [3:0] vns_videosoc_csrbank5_core_initiator_hres_backstore = 4'd0;
wire vns_videosoc_csrbank5_core_initiator_hres1_re;
wire [3:0] vns_videosoc_csrbank5_core_initiator_hres1_r;
wire [3:0] vns_videosoc_csrbank5_core_initiator_hres1_w;
wire vns_videosoc_csrbank5_core_initiator_hres0_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_hres0_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_hres0_w;
reg [3:0] vns_videosoc_csrbank5_core_initiator_hsync_start_backstore = 4'd0;
wire vns_videosoc_csrbank5_core_initiator_hsync_start1_re;
wire [3:0] vns_videosoc_csrbank5_core_initiator_hsync_start1_r;
wire [3:0] vns_videosoc_csrbank5_core_initiator_hsync_start1_w;
wire vns_videosoc_csrbank5_core_initiator_hsync_start0_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_hsync_start0_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_hsync_start0_w;
reg [3:0] vns_videosoc_csrbank5_core_initiator_hsync_end_backstore = 4'd0;
wire vns_videosoc_csrbank5_core_initiator_hsync_end1_re;
wire [3:0] vns_videosoc_csrbank5_core_initiator_hsync_end1_r;
wire [3:0] vns_videosoc_csrbank5_core_initiator_hsync_end1_w;
wire vns_videosoc_csrbank5_core_initiator_hsync_end0_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_hsync_end0_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_hsync_end0_w;
reg [3:0] vns_videosoc_csrbank5_core_initiator_hscan_backstore = 4'd0;
wire vns_videosoc_csrbank5_core_initiator_hscan1_re;
wire [3:0] vns_videosoc_csrbank5_core_initiator_hscan1_r;
wire [3:0] vns_videosoc_csrbank5_core_initiator_hscan1_w;
wire vns_videosoc_csrbank5_core_initiator_hscan0_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_hscan0_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_hscan0_w;
reg [3:0] vns_videosoc_csrbank5_core_initiator_vres_backstore = 4'd0;
wire vns_videosoc_csrbank5_core_initiator_vres1_re;
wire [3:0] vns_videosoc_csrbank5_core_initiator_vres1_r;
wire [3:0] vns_videosoc_csrbank5_core_initiator_vres1_w;
wire vns_videosoc_csrbank5_core_initiator_vres0_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_vres0_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_vres0_w;
reg [3:0] vns_videosoc_csrbank5_core_initiator_vsync_start_backstore = 4'd0;
wire vns_videosoc_csrbank5_core_initiator_vsync_start1_re;
wire [3:0] vns_videosoc_csrbank5_core_initiator_vsync_start1_r;
wire [3:0] vns_videosoc_csrbank5_core_initiator_vsync_start1_w;
wire vns_videosoc_csrbank5_core_initiator_vsync_start0_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_vsync_start0_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_vsync_start0_w;
reg [3:0] vns_videosoc_csrbank5_core_initiator_vsync_end_backstore = 4'd0;
wire vns_videosoc_csrbank5_core_initiator_vsync_end1_re;
wire [3:0] vns_videosoc_csrbank5_core_initiator_vsync_end1_r;
wire [3:0] vns_videosoc_csrbank5_core_initiator_vsync_end1_w;
wire vns_videosoc_csrbank5_core_initiator_vsync_end0_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_vsync_end0_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_vsync_end0_w;
reg [3:0] vns_videosoc_csrbank5_core_initiator_vscan_backstore = 4'd0;
wire vns_videosoc_csrbank5_core_initiator_vscan1_re;
wire [3:0] vns_videosoc_csrbank5_core_initiator_vscan1_r;
wire [3:0] vns_videosoc_csrbank5_core_initiator_vscan1_w;
wire vns_videosoc_csrbank5_core_initiator_vscan0_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_vscan0_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_vscan0_w;
reg [23:0] vns_videosoc_csrbank5_core_initiator_base_backstore = 24'd0;
wire vns_videosoc_csrbank5_core_initiator_base3_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_base3_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_base3_w;
wire vns_videosoc_csrbank5_core_initiator_base2_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_base2_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_base2_w;
wire vns_videosoc_csrbank5_core_initiator_base1_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_base1_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_base1_w;
wire vns_videosoc_csrbank5_core_initiator_base0_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_base0_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_base0_w;
reg [23:0] vns_videosoc_csrbank5_core_initiator_length_backstore = 24'd0;
wire vns_videosoc_csrbank5_core_initiator_length3_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_length3_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_length3_w;
wire vns_videosoc_csrbank5_core_initiator_length2_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_length2_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_length2_w;
wire vns_videosoc_csrbank5_core_initiator_length1_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_length1_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_length1_w;
wire vns_videosoc_csrbank5_core_initiator_length0_re;
wire [7:0] vns_videosoc_csrbank5_core_initiator_length0_r;
wire [7:0] vns_videosoc_csrbank5_core_initiator_length0_w;
wire vns_videosoc_csrbank5_driver_clocking_mmcm_reset0_re;
wire vns_videosoc_csrbank5_driver_clocking_mmcm_reset0_r;
wire vns_videosoc_csrbank5_driver_clocking_mmcm_reset0_w;
wire vns_videosoc_csrbank5_driver_clocking_mmcm_drdy_re;
wire vns_videosoc_csrbank5_driver_clocking_mmcm_drdy_r;
wire vns_videosoc_csrbank5_driver_clocking_mmcm_drdy_w;
wire vns_videosoc_csrbank5_driver_clocking_mmcm_adr0_re;
wire [6:0] vns_videosoc_csrbank5_driver_clocking_mmcm_adr0_r;
wire [6:0] vns_videosoc_csrbank5_driver_clocking_mmcm_adr0_w;
wire vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w1_re;
wire [7:0] vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w1_r;
wire [7:0] vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w1_w;
wire vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w0_re;
wire [7:0] vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w0_r;
wire [7:0] vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w0_w;
wire vns_videosoc_csrbank5_driver_clocking_mmcm_dat_r1_re;
wire [7:0] vns_videosoc_csrbank5_driver_clocking_mmcm_dat_r1_r;
wire [7:0] vns_videosoc_csrbank5_driver_clocking_mmcm_dat_r1_w;
wire vns_videosoc_csrbank5_driver_clocking_mmcm_dat_r0_re;
wire [7:0] vns_videosoc_csrbank5_driver_clocking_mmcm_dat_r0_r;
wire [7:0] vns_videosoc_csrbank5_driver_clocking_mmcm_dat_r0_w;
wire vns_videosoc_csrbank5_sel;
wire [13:0] vns_videosoc_interface6_bank_bus_adr;
wire vns_videosoc_interface6_bank_bus_we;
wire [7:0] vns_videosoc_interface6_bank_bus_dat_w;
reg [7:0] vns_videosoc_interface6_bank_bus_dat_r = 8'd0;
wire vns_videosoc_csrbank6_dna_id7_re;
wire vns_videosoc_csrbank6_dna_id7_r;
wire vns_videosoc_csrbank6_dna_id7_w;
wire vns_videosoc_csrbank6_dna_id6_re;
wire [7:0] vns_videosoc_csrbank6_dna_id6_r;
wire [7:0] vns_videosoc_csrbank6_dna_id6_w;
wire vns_videosoc_csrbank6_dna_id5_re;
wire [7:0] vns_videosoc_csrbank6_dna_id5_r;
wire [7:0] vns_videosoc_csrbank6_dna_id5_w;
wire vns_videosoc_csrbank6_dna_id4_re;
wire [7:0] vns_videosoc_csrbank6_dna_id4_r;
wire [7:0] vns_videosoc_csrbank6_dna_id4_w;
wire vns_videosoc_csrbank6_dna_id3_re;
wire [7:0] vns_videosoc_csrbank6_dna_id3_r;
wire [7:0] vns_videosoc_csrbank6_dna_id3_w;
wire vns_videosoc_csrbank6_dna_id2_re;
wire [7:0] vns_videosoc_csrbank6_dna_id2_r;
wire [7:0] vns_videosoc_csrbank6_dna_id2_w;
wire vns_videosoc_csrbank6_dna_id1_re;
wire [7:0] vns_videosoc_csrbank6_dna_id1_r;
wire [7:0] vns_videosoc_csrbank6_dna_id1_w;
wire vns_videosoc_csrbank6_dna_id0_re;
wire [7:0] vns_videosoc_csrbank6_dna_id0_r;
wire [7:0] vns_videosoc_csrbank6_dna_id0_w;
wire vns_videosoc_csrbank6_git_commit19_re;
wire [7:0] vns_videosoc_csrbank6_git_commit19_r;
wire [7:0] vns_videosoc_csrbank6_git_commit19_w;
wire vns_videosoc_csrbank6_git_commit18_re;
wire [7:0] vns_videosoc_csrbank6_git_commit18_r;
wire [7:0] vns_videosoc_csrbank6_git_commit18_w;
wire vns_videosoc_csrbank6_git_commit17_re;
wire [7:0] vns_videosoc_csrbank6_git_commit17_r;
wire [7:0] vns_videosoc_csrbank6_git_commit17_w;
wire vns_videosoc_csrbank6_git_commit16_re;
wire [7:0] vns_videosoc_csrbank6_git_commit16_r;
wire [7:0] vns_videosoc_csrbank6_git_commit16_w;
wire vns_videosoc_csrbank6_git_commit15_re;
wire [7:0] vns_videosoc_csrbank6_git_commit15_r;
wire [7:0] vns_videosoc_csrbank6_git_commit15_w;
wire vns_videosoc_csrbank6_git_commit14_re;
wire [7:0] vns_videosoc_csrbank6_git_commit14_r;
wire [7:0] vns_videosoc_csrbank6_git_commit14_w;
wire vns_videosoc_csrbank6_git_commit13_re;
wire [7:0] vns_videosoc_csrbank6_git_commit13_r;
wire [7:0] vns_videosoc_csrbank6_git_commit13_w;
wire vns_videosoc_csrbank6_git_commit12_re;
wire [7:0] vns_videosoc_csrbank6_git_commit12_r;
wire [7:0] vns_videosoc_csrbank6_git_commit12_w;
wire vns_videosoc_csrbank6_git_commit11_re;
wire [7:0] vns_videosoc_csrbank6_git_commit11_r;
wire [7:0] vns_videosoc_csrbank6_git_commit11_w;
wire vns_videosoc_csrbank6_git_commit10_re;
wire [7:0] vns_videosoc_csrbank6_git_commit10_r;
wire [7:0] vns_videosoc_csrbank6_git_commit10_w;
wire vns_videosoc_csrbank6_git_commit9_re;
wire [7:0] vns_videosoc_csrbank6_git_commit9_r;
wire [7:0] vns_videosoc_csrbank6_git_commit9_w;
wire vns_videosoc_csrbank6_git_commit8_re;
wire [7:0] vns_videosoc_csrbank6_git_commit8_r;
wire [7:0] vns_videosoc_csrbank6_git_commit8_w;
wire vns_videosoc_csrbank6_git_commit7_re;
wire [7:0] vns_videosoc_csrbank6_git_commit7_r;
wire [7:0] vns_videosoc_csrbank6_git_commit7_w;
wire vns_videosoc_csrbank6_git_commit6_re;
wire [7:0] vns_videosoc_csrbank6_git_commit6_r;
wire [7:0] vns_videosoc_csrbank6_git_commit6_w;
wire vns_videosoc_csrbank6_git_commit5_re;
wire [7:0] vns_videosoc_csrbank6_git_commit5_r;
wire [7:0] vns_videosoc_csrbank6_git_commit5_w;
wire vns_videosoc_csrbank6_git_commit4_re;
wire [7:0] vns_videosoc_csrbank6_git_commit4_r;
wire [7:0] vns_videosoc_csrbank6_git_commit4_w;
wire vns_videosoc_csrbank6_git_commit3_re;
wire [7:0] vns_videosoc_csrbank6_git_commit3_r;
wire [7:0] vns_videosoc_csrbank6_git_commit3_w;
wire vns_videosoc_csrbank6_git_commit2_re;
wire [7:0] vns_videosoc_csrbank6_git_commit2_r;
wire [7:0] vns_videosoc_csrbank6_git_commit2_w;
wire vns_videosoc_csrbank6_git_commit1_re;
wire [7:0] vns_videosoc_csrbank6_git_commit1_r;
wire [7:0] vns_videosoc_csrbank6_git_commit1_w;
wire vns_videosoc_csrbank6_git_commit0_re;
wire [7:0] vns_videosoc_csrbank6_git_commit0_r;
wire [7:0] vns_videosoc_csrbank6_git_commit0_w;
wire vns_videosoc_csrbank6_platform_platform7_re;
wire [7:0] vns_videosoc_csrbank6_platform_platform7_r;
wire [7:0] vns_videosoc_csrbank6_platform_platform7_w;
wire vns_videosoc_csrbank6_platform_platform6_re;
wire [7:0] vns_videosoc_csrbank6_platform_platform6_r;
wire [7:0] vns_videosoc_csrbank6_platform_platform6_w;
wire vns_videosoc_csrbank6_platform_platform5_re;
wire [7:0] vns_videosoc_csrbank6_platform_platform5_r;
wire [7:0] vns_videosoc_csrbank6_platform_platform5_w;
wire vns_videosoc_csrbank6_platform_platform4_re;
wire [7:0] vns_videosoc_csrbank6_platform_platform4_r;
wire [7:0] vns_videosoc_csrbank6_platform_platform4_w;
wire vns_videosoc_csrbank6_platform_platform3_re;
wire [7:0] vns_videosoc_csrbank6_platform_platform3_r;
wire [7:0] vns_videosoc_csrbank6_platform_platform3_w;
wire vns_videosoc_csrbank6_platform_platform2_re;
wire [7:0] vns_videosoc_csrbank6_platform_platform2_r;
wire [7:0] vns_videosoc_csrbank6_platform_platform2_w;
wire vns_videosoc_csrbank6_platform_platform1_re;
wire [7:0] vns_videosoc_csrbank6_platform_platform1_r;
wire [7:0] vns_videosoc_csrbank6_platform_platform1_w;
wire vns_videosoc_csrbank6_platform_platform0_re;
wire [7:0] vns_videosoc_csrbank6_platform_platform0_r;
wire [7:0] vns_videosoc_csrbank6_platform_platform0_w;
wire vns_videosoc_csrbank6_platform_target7_re;
wire [7:0] vns_videosoc_csrbank6_platform_target7_r;
wire [7:0] vns_videosoc_csrbank6_platform_target7_w;
wire vns_videosoc_csrbank6_platform_target6_re;
wire [7:0] vns_videosoc_csrbank6_platform_target6_r;
wire [7:0] vns_videosoc_csrbank6_platform_target6_w;
wire vns_videosoc_csrbank6_platform_target5_re;
wire [7:0] vns_videosoc_csrbank6_platform_target5_r;
wire [7:0] vns_videosoc_csrbank6_platform_target5_w;
wire vns_videosoc_csrbank6_platform_target4_re;
wire [7:0] vns_videosoc_csrbank6_platform_target4_r;
wire [7:0] vns_videosoc_csrbank6_platform_target4_w;
wire vns_videosoc_csrbank6_platform_target3_re;
wire [7:0] vns_videosoc_csrbank6_platform_target3_r;
wire [7:0] vns_videosoc_csrbank6_platform_target3_w;
wire vns_videosoc_csrbank6_platform_target2_re;
wire [7:0] vns_videosoc_csrbank6_platform_target2_r;
wire [7:0] vns_videosoc_csrbank6_platform_target2_w;
wire vns_videosoc_csrbank6_platform_target1_re;
wire [7:0] vns_videosoc_csrbank6_platform_target1_r;
wire [7:0] vns_videosoc_csrbank6_platform_target1_w;
wire vns_videosoc_csrbank6_platform_target0_re;
wire [7:0] vns_videosoc_csrbank6_platform_target0_r;
wire [7:0] vns_videosoc_csrbank6_platform_target0_w;
wire vns_videosoc_csrbank6_xadc_temperature1_re;
wire [3:0] vns_videosoc_csrbank6_xadc_temperature1_r;
wire [3:0] vns_videosoc_csrbank6_xadc_temperature1_w;
wire vns_videosoc_csrbank6_xadc_temperature0_re;
wire [7:0] vns_videosoc_csrbank6_xadc_temperature0_r;
wire [7:0] vns_videosoc_csrbank6_xadc_temperature0_w;
wire vns_videosoc_csrbank6_xadc_vccint1_re;
wire [3:0] vns_videosoc_csrbank6_xadc_vccint1_r;
wire [3:0] vns_videosoc_csrbank6_xadc_vccint1_w;
wire vns_videosoc_csrbank6_xadc_vccint0_re;
wire [7:0] vns_videosoc_csrbank6_xadc_vccint0_r;
wire [7:0] vns_videosoc_csrbank6_xadc_vccint0_w;
wire vns_videosoc_csrbank6_xadc_vccaux1_re;
wire [3:0] vns_videosoc_csrbank6_xadc_vccaux1_r;
wire [3:0] vns_videosoc_csrbank6_xadc_vccaux1_w;
wire vns_videosoc_csrbank6_xadc_vccaux0_re;
wire [7:0] vns_videosoc_csrbank6_xadc_vccaux0_r;
wire [7:0] vns_videosoc_csrbank6_xadc_vccaux0_w;
wire vns_videosoc_csrbank6_xadc_vccbram1_re;
wire [3:0] vns_videosoc_csrbank6_xadc_vccbram1_r;
wire [3:0] vns_videosoc_csrbank6_xadc_vccbram1_w;
wire vns_videosoc_csrbank6_xadc_vccbram0_re;
wire [7:0] vns_videosoc_csrbank6_xadc_vccbram0_r;
wire [7:0] vns_videosoc_csrbank6_xadc_vccbram0_w;
wire vns_videosoc_csrbank6_sel;
wire [13:0] vns_videosoc_interface7_bank_bus_adr;
wire vns_videosoc_interface7_bank_bus_we;
wire [7:0] vns_videosoc_interface7_bank_bus_dat_w;
reg [7:0] vns_videosoc_interface7_bank_bus_dat_r = 8'd0;
wire vns_videosoc_csrbank7_spi_length0_re;
wire [7:0] vns_videosoc_csrbank7_spi_length0_r;
wire [7:0] vns_videosoc_csrbank7_spi_length0_w;
wire vns_videosoc_csrbank7_spi_status_re;
wire vns_videosoc_csrbank7_spi_status_r;
wire vns_videosoc_csrbank7_spi_status_w;
wire vns_videosoc_csrbank7_spi_mosi0_re;
wire [7:0] vns_videosoc_csrbank7_spi_mosi0_r;
wire [7:0] vns_videosoc_csrbank7_spi_mosi0_w;
wire vns_videosoc_csrbank7_gpio_out0_re;
wire [3:0] vns_videosoc_csrbank7_gpio_out0_r;
wire [3:0] vns_videosoc_csrbank7_gpio_out0_w;
wire vns_videosoc_csrbank7_sel;
wire [13:0] vns_videosoc_interface8_bank_bus_adr;
wire vns_videosoc_interface8_bank_bus_we;
wire [7:0] vns_videosoc_interface8_bank_bus_dat_w;
reg [7:0] vns_videosoc_interface8_bank_bus_dat_r = 8'd0;
wire vns_videosoc_csrbank8_dfii_control0_re;
wire [3:0] vns_videosoc_csrbank8_dfii_control0_r;
wire [3:0] vns_videosoc_csrbank8_dfii_control0_w;
wire vns_videosoc_csrbank8_dfii_pi0_command0_re;
wire [5:0] vns_videosoc_csrbank8_dfii_pi0_command0_r;
wire [5:0] vns_videosoc_csrbank8_dfii_pi0_command0_w;
wire vns_videosoc_csrbank8_dfii_pi0_address1_re;
wire [6:0] vns_videosoc_csrbank8_dfii_pi0_address1_r;
wire [6:0] vns_videosoc_csrbank8_dfii_pi0_address1_w;
wire vns_videosoc_csrbank8_dfii_pi0_address0_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_address0_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_address0_w;
wire vns_videosoc_csrbank8_dfii_pi0_baddress0_re;
wire [2:0] vns_videosoc_csrbank8_dfii_pi0_baddress0_r;
wire [2:0] vns_videosoc_csrbank8_dfii_pi0_baddress0_w;
wire vns_videosoc_csrbank8_dfii_pi0_wrdata3_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_wrdata3_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_wrdata3_w;
wire vns_videosoc_csrbank8_dfii_pi0_wrdata2_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_wrdata2_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_wrdata2_w;
wire vns_videosoc_csrbank8_dfii_pi0_wrdata1_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_wrdata1_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_wrdata1_w;
wire vns_videosoc_csrbank8_dfii_pi0_wrdata0_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_wrdata0_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_wrdata0_w;
wire vns_videosoc_csrbank8_dfii_pi0_rddata3_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_rddata3_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_rddata3_w;
wire vns_videosoc_csrbank8_dfii_pi0_rddata2_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_rddata2_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_rddata2_w;
wire vns_videosoc_csrbank8_dfii_pi0_rddata1_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_rddata1_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_rddata1_w;
wire vns_videosoc_csrbank8_dfii_pi0_rddata0_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_rddata0_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi0_rddata0_w;
wire vns_videosoc_csrbank8_dfii_pi1_command0_re;
wire [5:0] vns_videosoc_csrbank8_dfii_pi1_command0_r;
wire [5:0] vns_videosoc_csrbank8_dfii_pi1_command0_w;
wire vns_videosoc_csrbank8_dfii_pi1_address1_re;
wire [6:0] vns_videosoc_csrbank8_dfii_pi1_address1_r;
wire [6:0] vns_videosoc_csrbank8_dfii_pi1_address1_w;
wire vns_videosoc_csrbank8_dfii_pi1_address0_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_address0_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_address0_w;
wire vns_videosoc_csrbank8_dfii_pi1_baddress0_re;
wire [2:0] vns_videosoc_csrbank8_dfii_pi1_baddress0_r;
wire [2:0] vns_videosoc_csrbank8_dfii_pi1_baddress0_w;
wire vns_videosoc_csrbank8_dfii_pi1_wrdata3_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_wrdata3_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_wrdata3_w;
wire vns_videosoc_csrbank8_dfii_pi1_wrdata2_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_wrdata2_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_wrdata2_w;
wire vns_videosoc_csrbank8_dfii_pi1_wrdata1_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_wrdata1_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_wrdata1_w;
wire vns_videosoc_csrbank8_dfii_pi1_wrdata0_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_wrdata0_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_wrdata0_w;
wire vns_videosoc_csrbank8_dfii_pi1_rddata3_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_rddata3_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_rddata3_w;
wire vns_videosoc_csrbank8_dfii_pi1_rddata2_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_rddata2_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_rddata2_w;
wire vns_videosoc_csrbank8_dfii_pi1_rddata1_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_rddata1_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_rddata1_w;
wire vns_videosoc_csrbank8_dfii_pi1_rddata0_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_rddata0_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi1_rddata0_w;
wire vns_videosoc_csrbank8_dfii_pi2_command0_re;
wire [5:0] vns_videosoc_csrbank8_dfii_pi2_command0_r;
wire [5:0] vns_videosoc_csrbank8_dfii_pi2_command0_w;
wire vns_videosoc_csrbank8_dfii_pi2_address1_re;
wire [6:0] vns_videosoc_csrbank8_dfii_pi2_address1_r;
wire [6:0] vns_videosoc_csrbank8_dfii_pi2_address1_w;
wire vns_videosoc_csrbank8_dfii_pi2_address0_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_address0_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_address0_w;
wire vns_videosoc_csrbank8_dfii_pi2_baddress0_re;
wire [2:0] vns_videosoc_csrbank8_dfii_pi2_baddress0_r;
wire [2:0] vns_videosoc_csrbank8_dfii_pi2_baddress0_w;
wire vns_videosoc_csrbank8_dfii_pi2_wrdata3_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_wrdata3_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_wrdata3_w;
wire vns_videosoc_csrbank8_dfii_pi2_wrdata2_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_wrdata2_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_wrdata2_w;
wire vns_videosoc_csrbank8_dfii_pi2_wrdata1_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_wrdata1_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_wrdata1_w;
wire vns_videosoc_csrbank8_dfii_pi2_wrdata0_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_wrdata0_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_wrdata0_w;
wire vns_videosoc_csrbank8_dfii_pi2_rddata3_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_rddata3_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_rddata3_w;
wire vns_videosoc_csrbank8_dfii_pi2_rddata2_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_rddata2_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_rddata2_w;
wire vns_videosoc_csrbank8_dfii_pi2_rddata1_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_rddata1_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_rddata1_w;
wire vns_videosoc_csrbank8_dfii_pi2_rddata0_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_rddata0_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi2_rddata0_w;
wire vns_videosoc_csrbank8_dfii_pi3_command0_re;
wire [5:0] vns_videosoc_csrbank8_dfii_pi3_command0_r;
wire [5:0] vns_videosoc_csrbank8_dfii_pi3_command0_w;
wire vns_videosoc_csrbank8_dfii_pi3_address1_re;
wire [6:0] vns_videosoc_csrbank8_dfii_pi3_address1_r;
wire [6:0] vns_videosoc_csrbank8_dfii_pi3_address1_w;
wire vns_videosoc_csrbank8_dfii_pi3_address0_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_address0_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_address0_w;
wire vns_videosoc_csrbank8_dfii_pi3_baddress0_re;
wire [2:0] vns_videosoc_csrbank8_dfii_pi3_baddress0_r;
wire [2:0] vns_videosoc_csrbank8_dfii_pi3_baddress0_w;
wire vns_videosoc_csrbank8_dfii_pi3_wrdata3_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_wrdata3_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_wrdata3_w;
wire vns_videosoc_csrbank8_dfii_pi3_wrdata2_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_wrdata2_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_wrdata2_w;
wire vns_videosoc_csrbank8_dfii_pi3_wrdata1_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_wrdata1_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_wrdata1_w;
wire vns_videosoc_csrbank8_dfii_pi3_wrdata0_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_wrdata0_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_wrdata0_w;
wire vns_videosoc_csrbank8_dfii_pi3_rddata3_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_rddata3_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_rddata3_w;
wire vns_videosoc_csrbank8_dfii_pi3_rddata2_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_rddata2_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_rddata2_w;
wire vns_videosoc_csrbank8_dfii_pi3_rddata1_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_rddata1_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_rddata1_w;
wire vns_videosoc_csrbank8_dfii_pi3_rddata0_re;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_rddata0_r;
wire [7:0] vns_videosoc_csrbank8_dfii_pi3_rddata0_w;
wire vns_videosoc_csrbank8_controller_bandwidth_nreads2_re;
wire [7:0] vns_videosoc_csrbank8_controller_bandwidth_nreads2_r;
wire [7:0] vns_videosoc_csrbank8_controller_bandwidth_nreads2_w;
wire vns_videosoc_csrbank8_controller_bandwidth_nreads1_re;
wire [7:0] vns_videosoc_csrbank8_controller_bandwidth_nreads1_r;
wire [7:0] vns_videosoc_csrbank8_controller_bandwidth_nreads1_w;
wire vns_videosoc_csrbank8_controller_bandwidth_nreads0_re;
wire [7:0] vns_videosoc_csrbank8_controller_bandwidth_nreads0_r;
wire [7:0] vns_videosoc_csrbank8_controller_bandwidth_nreads0_w;
wire vns_videosoc_csrbank8_controller_bandwidth_nwrites2_re;
wire [7:0] vns_videosoc_csrbank8_controller_bandwidth_nwrites2_r;
wire [7:0] vns_videosoc_csrbank8_controller_bandwidth_nwrites2_w;
wire vns_videosoc_csrbank8_controller_bandwidth_nwrites1_re;
wire [7:0] vns_videosoc_csrbank8_controller_bandwidth_nwrites1_r;
wire [7:0] vns_videosoc_csrbank8_controller_bandwidth_nwrites1_w;
wire vns_videosoc_csrbank8_controller_bandwidth_nwrites0_re;
wire [7:0] vns_videosoc_csrbank8_controller_bandwidth_nwrites0_r;
wire [7:0] vns_videosoc_csrbank8_controller_bandwidth_nwrites0_w;
wire vns_videosoc_csrbank8_controller_bandwidth_data_width_re;
wire [7:0] vns_videosoc_csrbank8_controller_bandwidth_data_width_r;
wire [7:0] vns_videosoc_csrbank8_controller_bandwidth_data_width_w;
wire vns_videosoc_csrbank8_sel;
wire [13:0] vns_videosoc_interface9_bank_bus_adr;
wire vns_videosoc_interface9_bank_bus_we;
wire [7:0] vns_videosoc_interface9_bank_bus_dat_w;
reg [7:0] vns_videosoc_interface9_bank_bus_dat_r = 8'd0;
wire vns_videosoc_csrbank9_bitbang0_re;
wire [3:0] vns_videosoc_csrbank9_bitbang0_r;
wire [3:0] vns_videosoc_csrbank9_bitbang0_w;
wire vns_videosoc_csrbank9_miso_re;
wire vns_videosoc_csrbank9_miso_r;
wire vns_videosoc_csrbank9_miso_w;
wire vns_videosoc_csrbank9_bitbang_en0_re;
wire vns_videosoc_csrbank9_bitbang_en0_r;
wire vns_videosoc_csrbank9_bitbang_en0_w;
wire vns_videosoc_csrbank9_sel;
wire [13:0] vns_videosoc_interface10_bank_bus_adr;
wire vns_videosoc_interface10_bank_bus_we;
wire [7:0] vns_videosoc_interface10_bank_bus_dat_w;
reg [7:0] vns_videosoc_interface10_bank_bus_dat_r = 8'd0;
wire vns_videosoc_csrbank10_load3_re;
wire [7:0] vns_videosoc_csrbank10_load3_r;
wire [7:0] vns_videosoc_csrbank10_load3_w;
wire vns_videosoc_csrbank10_load2_re;
wire [7:0] vns_videosoc_csrbank10_load2_r;
wire [7:0] vns_videosoc_csrbank10_load2_w;
wire vns_videosoc_csrbank10_load1_re;
wire [7:0] vns_videosoc_csrbank10_load1_r;
wire [7:0] vns_videosoc_csrbank10_load1_w;
wire vns_videosoc_csrbank10_load0_re;
wire [7:0] vns_videosoc_csrbank10_load0_r;
wire [7:0] vns_videosoc_csrbank10_load0_w;
wire vns_videosoc_csrbank10_reload3_re;
wire [7:0] vns_videosoc_csrbank10_reload3_r;
wire [7:0] vns_videosoc_csrbank10_reload3_w;
wire vns_videosoc_csrbank10_reload2_re;
wire [7:0] vns_videosoc_csrbank10_reload2_r;
wire [7:0] vns_videosoc_csrbank10_reload2_w;
wire vns_videosoc_csrbank10_reload1_re;
wire [7:0] vns_videosoc_csrbank10_reload1_r;
wire [7:0] vns_videosoc_csrbank10_reload1_w;
wire vns_videosoc_csrbank10_reload0_re;
wire [7:0] vns_videosoc_csrbank10_reload0_r;
wire [7:0] vns_videosoc_csrbank10_reload0_w;
wire vns_videosoc_csrbank10_en0_re;
wire vns_videosoc_csrbank10_en0_r;
wire vns_videosoc_csrbank10_en0_w;
wire vns_videosoc_csrbank10_value3_re;
wire [7:0] vns_videosoc_csrbank10_value3_r;
wire [7:0] vns_videosoc_csrbank10_value3_w;
wire vns_videosoc_csrbank10_value2_re;
wire [7:0] vns_videosoc_csrbank10_value2_r;
wire [7:0] vns_videosoc_csrbank10_value2_w;
wire vns_videosoc_csrbank10_value1_re;
wire [7:0] vns_videosoc_csrbank10_value1_r;
wire [7:0] vns_videosoc_csrbank10_value1_w;
wire vns_videosoc_csrbank10_value0_re;
wire [7:0] vns_videosoc_csrbank10_value0_r;
wire [7:0] vns_videosoc_csrbank10_value0_w;
wire vns_videosoc_csrbank10_ev_enable0_re;
wire vns_videosoc_csrbank10_ev_enable0_r;
wire vns_videosoc_csrbank10_ev_enable0_w;
wire vns_videosoc_csrbank10_sel;
wire [13:0] vns_videosoc_interface11_bank_bus_adr;
wire vns_videosoc_interface11_bank_bus_we;
wire [7:0] vns_videosoc_interface11_bank_bus_dat_w;
reg [7:0] vns_videosoc_interface11_bank_bus_dat_r = 8'd0;
wire vns_videosoc_csrbank11_txfull_re;
wire vns_videosoc_csrbank11_txfull_r;
wire vns_videosoc_csrbank11_txfull_w;
wire vns_videosoc_csrbank11_rxempty_re;
wire vns_videosoc_csrbank11_rxempty_r;
wire vns_videosoc_csrbank11_rxempty_w;
wire vns_videosoc_csrbank11_ev_enable0_re;
wire [1:0] vns_videosoc_csrbank11_ev_enable0_r;
wire [1:0] vns_videosoc_csrbank11_ev_enable0_w;
wire vns_videosoc_csrbank11_sel;
wire [13:0] vns_videosoc_interface12_bank_bus_adr;
wire vns_videosoc_interface12_bank_bus_we;
wire [7:0] vns_videosoc_interface12_bank_bus_dat_w;
reg [7:0] vns_videosoc_interface12_bank_bus_dat_r = 8'd0;
wire vns_videosoc_csrbank12_tuning_word3_re;
wire [7:0] vns_videosoc_csrbank12_tuning_word3_r;
wire [7:0] vns_videosoc_csrbank12_tuning_word3_w;
wire vns_videosoc_csrbank12_tuning_word2_re;
wire [7:0] vns_videosoc_csrbank12_tuning_word2_r;
wire [7:0] vns_videosoc_csrbank12_tuning_word2_w;
wire vns_videosoc_csrbank12_tuning_word1_re;
wire [7:0] vns_videosoc_csrbank12_tuning_word1_r;
wire [7:0] vns_videosoc_csrbank12_tuning_word1_w;
wire vns_videosoc_csrbank12_tuning_word0_re;
wire [7:0] vns_videosoc_csrbank12_tuning_word0_r;
wire [7:0] vns_videosoc_csrbank12_tuning_word0_w;
wire vns_videosoc_csrbank12_sel;
reg vns_comb_rhs_array_muxed0 = 1'd0;
reg [14:0] vns_comb_rhs_array_muxed1 = 15'd0;
reg [2:0] vns_comb_rhs_array_muxed2 = 3'd0;
reg vns_comb_rhs_array_muxed3 = 1'd0;
reg vns_comb_rhs_array_muxed4 = 1'd0;
reg vns_comb_rhs_array_muxed5 = 1'd0;
reg vns_comb_t_array_muxed0 = 1'd0;
reg vns_comb_t_array_muxed1 = 1'd0;
reg vns_comb_t_array_muxed2 = 1'd0;
reg vns_comb_rhs_array_muxed6 = 1'd0;
reg [14:0] vns_comb_rhs_array_muxed7 = 15'd0;
reg [2:0] vns_comb_rhs_array_muxed8 = 3'd0;
reg vns_comb_rhs_array_muxed9 = 1'd0;
reg vns_comb_rhs_array_muxed10 = 1'd0;
reg vns_comb_rhs_array_muxed11 = 1'd0;
reg vns_comb_t_array_muxed3 = 1'd0;
reg vns_comb_t_array_muxed4 = 1'd0;
reg vns_comb_t_array_muxed5 = 1'd0;
reg [21:0] vns_comb_rhs_array_muxed12 = 22'd0;
reg vns_comb_rhs_array_muxed13 = 1'd0;
reg vns_comb_rhs_array_muxed14 = 1'd0;
reg [21:0] vns_comb_rhs_array_muxed15 = 22'd0;
reg vns_comb_rhs_array_muxed16 = 1'd0;
reg vns_comb_rhs_array_muxed17 = 1'd0;
reg [21:0] vns_comb_rhs_array_muxed18 = 22'd0;
reg vns_comb_rhs_array_muxed19 = 1'd0;
reg vns_comb_rhs_array_muxed20 = 1'd0;
reg [21:0] vns_comb_rhs_array_muxed21 = 22'd0;
reg vns_comb_rhs_array_muxed22 = 1'd0;
reg vns_comb_rhs_array_muxed23 = 1'd0;
reg [21:0] vns_comb_rhs_array_muxed24 = 22'd0;
reg vns_comb_rhs_array_muxed25 = 1'd0;
reg vns_comb_rhs_array_muxed26 = 1'd0;
reg [21:0] vns_comb_rhs_array_muxed27 = 22'd0;
reg vns_comb_rhs_array_muxed28 = 1'd0;
reg vns_comb_rhs_array_muxed29 = 1'd0;
reg [21:0] vns_comb_rhs_array_muxed30 = 22'd0;
reg vns_comb_rhs_array_muxed31 = 1'd0;
reg vns_comb_rhs_array_muxed32 = 1'd0;
reg [21:0] vns_comb_rhs_array_muxed33 = 22'd0;
reg vns_comb_rhs_array_muxed34 = 1'd0;
reg vns_comb_rhs_array_muxed35 = 1'd0;
reg [24:0] vns_comb_rhs_array_muxed36 = 25'd0;
reg vns_comb_rhs_array_muxed37 = 1'd0;
reg [29:0] vns_comb_rhs_array_muxed38 = 30'd0;
reg [31:0] vns_comb_rhs_array_muxed39 = 32'd0;
reg [3:0] vns_comb_rhs_array_muxed40 = 4'd0;
reg vns_comb_rhs_array_muxed41 = 1'd0;
reg vns_comb_rhs_array_muxed42 = 1'd0;
reg vns_comb_rhs_array_muxed43 = 1'd0;
reg [2:0] vns_comb_rhs_array_muxed44 = 3'd0;
reg [1:0] vns_comb_rhs_array_muxed45 = 2'd0;
reg [29:0] vns_comb_rhs_array_muxed46 = 30'd0;
reg [31:0] vns_comb_rhs_array_muxed47 = 32'd0;
reg [3:0] vns_comb_rhs_array_muxed48 = 4'd0;
reg vns_comb_rhs_array_muxed49 = 1'd0;
reg vns_comb_rhs_array_muxed50 = 1'd0;
reg vns_comb_rhs_array_muxed51 = 1'd0;
reg [2:0] vns_comb_rhs_array_muxed52 = 3'd0;
reg [1:0] vns_comb_rhs_array_muxed53 = 2'd0;
reg [9:0] vns_sync_f_array_muxed0 = 10'd0;
reg [9:0] vns_sync_f_array_muxed1 = 10'd0;
reg [9:0] vns_sync_f_array_muxed2 = 10'd0;
reg [14:0] vns_sync_rhs_array_muxed0 = 15'd0;
reg [2:0] vns_sync_rhs_array_muxed1 = 3'd0;
reg vns_sync_rhs_array_muxed2 = 1'd0;
reg vns_sync_rhs_array_muxed3 = 1'd0;
reg vns_sync_rhs_array_muxed4 = 1'd0;
reg vns_sync_rhs_array_muxed5 = 1'd0;
reg vns_sync_rhs_array_muxed6 = 1'd0;
reg [14:0] vns_sync_rhs_array_muxed7 = 15'd0;
reg [2:0] vns_sync_rhs_array_muxed8 = 3'd0;
reg vns_sync_rhs_array_muxed9 = 1'd0;
reg vns_sync_rhs_array_muxed10 = 1'd0;
reg vns_sync_rhs_array_muxed11 = 1'd0;
reg vns_sync_rhs_array_muxed12 = 1'd0;
reg vns_sync_rhs_array_muxed13 = 1'd0;
reg [14:0] vns_sync_rhs_array_muxed14 = 15'd0;
reg [2:0] vns_sync_rhs_array_muxed15 = 3'd0;
reg vns_sync_rhs_array_muxed16 = 1'd0;
reg vns_sync_rhs_array_muxed17 = 1'd0;
reg vns_sync_rhs_array_muxed18 = 1'd0;
reg vns_sync_rhs_array_muxed19 = 1'd0;
reg vns_sync_rhs_array_muxed20 = 1'd0;
reg [14:0] vns_sync_rhs_array_muxed21 = 15'd0;
reg [2:0] vns_sync_rhs_array_muxed22 = 3'd0;
reg vns_sync_rhs_array_muxed23 = 1'd0;
reg vns_sync_rhs_array_muxed24 = 1'd0;
reg vns_sync_rhs_array_muxed25 = 1'd0;
reg vns_sync_rhs_array_muxed26 = 1'd0;
reg vns_sync_rhs_array_muxed27 = 1'd0;
(* ars_false_path = "true" *) wire vns_xilinxasyncresetsynchronizerimpl0;
wire vns_xilinxasyncresetsynchronizerimpl0_rst_meta;
(* ars_false_path = "true" *) wire vns_xilinxasyncresetsynchronizerimpl1;
wire vns_xilinxasyncresetsynchronizerimpl1_rst_meta;
(* ars_false_path = "true" *) wire vns_xilinxasyncresetsynchronizerimpl2;
wire vns_xilinxasyncresetsynchronizerimpl2_rst_meta;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl0_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl0_regs1 = 1'd0;
wire vns_xilinxasyncresetsynchronizerimpl3_rst_meta;
wire vns_xilinxasyncresetsynchronizerimpl4_rst_meta;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl1_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl1_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl2_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl2_regs1 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl3_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl3_regs1 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl4_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl4_regs1 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl5_regs0 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg [6:0] vns_xilinxmultiregimpl5_regs1 = 7'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl6_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl6_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl7_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl7_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl8_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl8_regs1 = 1'd0;
(* ars_false_path = "true" *) wire vns_xilinxasyncresetsynchronizerimpl5;
wire vns_xilinxasyncresetsynchronizerimpl5_rst_meta;
(* ars_false_path = "true" *) wire vns_xilinxasyncresetsynchronizerimpl6;
wire vns_xilinxasyncresetsynchronizerimpl6_rst_meta;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl9_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl9_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl10_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl10_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl11_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl11_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl12_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl12_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl13_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl13_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl14_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl14_regs1 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl15_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl15_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl16_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl16_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl17_regs0 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl17_regs1 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl18_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl18_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl19_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl19_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl20_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl20_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl21_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl21_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl22_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl22_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl23_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl23_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl24_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl24_regs1 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl25_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl25_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl26_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl26_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl27_regs0 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl27_regs1 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl28_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl28_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl29_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl29_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl30_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl30_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl31_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl31_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl32_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl32_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl33_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl33_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl34_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl34_regs1 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl35_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl35_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl36_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl36_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl37_regs0 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg [3:0] vns_xilinxmultiregimpl37_regs1 = 4'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl38_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl38_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl39_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl39_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl40_regs0 = 11'd0;
(* async_reg = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl40_regs1 = 11'd0;
(* async_reg = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl41_regs0 = 11'd0;
(* async_reg = "true", dont_touch = "true" *) reg [10:0] vns_xilinxmultiregimpl41_regs1 = 11'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] vns_xilinxmultiregimpl42_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] vns_xilinxmultiregimpl42_regs1 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] vns_xilinxmultiregimpl43_regs0 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg [9:0] vns_xilinxmultiregimpl43_regs1 = 10'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl44_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl44_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl45_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl45_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl46_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl46_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg [5:0] vns_xilinxmultiregimpl47_regs0 = 6'd0;
(* async_reg = "true", dont_touch = "true" *) reg [5:0] vns_xilinxmultiregimpl47_regs1 = 6'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl48_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl48_regs1 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl49_regs0 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [2:0] vns_xilinxmultiregimpl49_regs1 = 3'd0;
(* async_reg = "true", dont_touch = "true" *) reg [4:0] vns_xilinxmultiregimpl50_regs0 = 5'd0;
(* async_reg = "true", dont_touch = "true" *) reg [4:0] vns_xilinxmultiregimpl50_regs1 = 5'd0;
(* async_reg = "true", dont_touch = "true" *) reg [4:0] vns_xilinxmultiregimpl51_regs0 = 5'd0;
(* async_reg = "true", dont_touch = "true" *) reg [4:0] vns_xilinxmultiregimpl51_regs1 = 5'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl52_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl52_regs1 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl53_regs0 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg [1:0] vns_xilinxmultiregimpl53_regs1 = 2'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl54_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl54_regs1 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl55_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg vns_xilinxmultiregimpl55_regs1 = 1'd0;

assign soc_videosoc_sel = user_sw0;
assign soc_hdmi_in0_freq_clk0 = hdmi_in0_pix_clk;
assign hdmi_in_txen = 1'd1;
always @(*) begin
	soc_videosoc_videosoc_interrupt <= 32'd0;
	soc_videosoc_videosoc_interrupt[1] <= soc_videosoc_videosoc_irq;
	soc_videosoc_videosoc_interrupt[2] <= soc_videosoc_uart_irq;
	soc_videosoc_videosoc_interrupt[3] <= soc_ethmac_ev_irq;
	soc_videosoc_videosoc_interrupt[4] <= soc_dma_slot_array_irq;
end
assign soc_videosoc_videosoc_ibus_adr = soc_videosoc_videosoc_i_adr_o[31:2];
assign soc_videosoc_videosoc_dbus_adr = soc_videosoc_videosoc_d_adr_o[31:2];
assign soc_videosoc_videosoc_rom_adr = soc_videosoc_videosoc_rom_bus_adr[12:0];
assign soc_videosoc_videosoc_rom_bus_dat_r = soc_videosoc_videosoc_rom_dat_r;
always @(*) begin
	soc_videosoc_videosoc_sram_we <= 4'd0;
	soc_videosoc_videosoc_sram_we[0] <= (((soc_videosoc_videosoc_sram_bus_cyc & soc_videosoc_videosoc_sram_bus_stb) & soc_videosoc_videosoc_sram_bus_we) & soc_videosoc_videosoc_sram_bus_sel[0]);
	soc_videosoc_videosoc_sram_we[1] <= (((soc_videosoc_videosoc_sram_bus_cyc & soc_videosoc_videosoc_sram_bus_stb) & soc_videosoc_videosoc_sram_bus_we) & soc_videosoc_videosoc_sram_bus_sel[1]);
	soc_videosoc_videosoc_sram_we[2] <= (((soc_videosoc_videosoc_sram_bus_cyc & soc_videosoc_videosoc_sram_bus_stb) & soc_videosoc_videosoc_sram_bus_we) & soc_videosoc_videosoc_sram_bus_sel[2]);
	soc_videosoc_videosoc_sram_we[3] <= (((soc_videosoc_videosoc_sram_bus_cyc & soc_videosoc_videosoc_sram_bus_stb) & soc_videosoc_videosoc_sram_bus_we) & soc_videosoc_videosoc_sram_bus_sel[3]);
end
assign soc_videosoc_videosoc_sram_adr = soc_videosoc_videosoc_sram_bus_adr[12:0];
assign soc_videosoc_videosoc_sram_bus_dat_r = soc_videosoc_videosoc_sram_dat_r;
assign soc_videosoc_videosoc_sram_dat_w = soc_videosoc_videosoc_sram_bus_dat_w;
assign soc_videosoc_videosoc_zero_trigger = (soc_videosoc_videosoc_value != 1'd0);
assign soc_videosoc_videosoc_eventmanager_status_w = soc_videosoc_videosoc_zero_status;
always @(*) begin
	soc_videosoc_videosoc_zero_clear <= 1'd0;
	if ((soc_videosoc_videosoc_eventmanager_pending_re & soc_videosoc_videosoc_eventmanager_pending_r)) begin
		soc_videosoc_videosoc_zero_clear <= 1'd1;
	end
end
assign soc_videosoc_videosoc_eventmanager_pending_w = soc_videosoc_videosoc_zero_pending;
assign soc_videosoc_videosoc_irq = (soc_videosoc_videosoc_eventmanager_pending_w & soc_videosoc_videosoc_eventmanager_storage);
assign soc_videosoc_videosoc_zero_status = soc_videosoc_videosoc_zero_trigger;
assign soc_videosoc_uart_tx_fifo_sink_valid = soc_videosoc_uart_rxtx_re;
assign soc_videosoc_uart_tx_fifo_sink_payload_data = soc_videosoc_uart_rxtx_r;
assign soc_videosoc_uart_txfull_status = (~soc_videosoc_uart_tx_fifo_sink_ready);
assign soc_videosoc_rs232phyinterface0_sink_valid = soc_videosoc_uart_tx_fifo_source_valid;
assign soc_videosoc_uart_tx_fifo_source_ready = soc_videosoc_rs232phyinterface0_sink_ready;
assign soc_videosoc_rs232phyinterface0_sink_first = soc_videosoc_uart_tx_fifo_source_first;
assign soc_videosoc_rs232phyinterface0_sink_last = soc_videosoc_uart_tx_fifo_source_last;
assign soc_videosoc_rs232phyinterface0_sink_payload_data = soc_videosoc_uart_tx_fifo_source_payload_data;
assign soc_videosoc_uart_tx_trigger = (~soc_videosoc_uart_tx_fifo_sink_ready);
assign soc_videosoc_uart_rx_fifo_sink_valid = soc_videosoc_rs232phyinterface0_source_valid;
assign soc_videosoc_rs232phyinterface0_source_ready = soc_videosoc_uart_rx_fifo_sink_ready;
assign soc_videosoc_uart_rx_fifo_sink_first = soc_videosoc_rs232phyinterface0_source_first;
assign soc_videosoc_uart_rx_fifo_sink_last = soc_videosoc_rs232phyinterface0_source_last;
assign soc_videosoc_uart_rx_fifo_sink_payload_data = soc_videosoc_rs232phyinterface0_source_payload_data;
assign soc_videosoc_uart_rxempty_status = (~soc_videosoc_uart_rx_fifo_source_valid);
assign soc_videosoc_uart_rxtx_w = soc_videosoc_uart_rx_fifo_source_payload_data;
assign soc_videosoc_uart_rx_fifo_source_ready = soc_videosoc_uart_rx_clear;
assign soc_videosoc_uart_rx_trigger = (~soc_videosoc_uart_rx_fifo_source_valid);
always @(*) begin
	soc_videosoc_uart_tx_clear <= 1'd0;
	if ((soc_videosoc_uart_pending_re & soc_videosoc_uart_pending_r[0])) begin
		soc_videosoc_uart_tx_clear <= 1'd1;
	end
end
always @(*) begin
	soc_videosoc_uart_status_w <= 2'd0;
	soc_videosoc_uart_status_w[0] <= soc_videosoc_uart_tx_status;
	soc_videosoc_uart_status_w[1] <= soc_videosoc_uart_rx_status;
end
always @(*) begin
	soc_videosoc_uart_rx_clear <= 1'd0;
	if ((soc_videosoc_uart_pending_re & soc_videosoc_uart_pending_r[1])) begin
		soc_videosoc_uart_rx_clear <= 1'd1;
	end
end
always @(*) begin
	soc_videosoc_uart_pending_w <= 2'd0;
	soc_videosoc_uart_pending_w[0] <= soc_videosoc_uart_tx_pending;
	soc_videosoc_uart_pending_w[1] <= soc_videosoc_uart_rx_pending;
end
assign soc_videosoc_uart_irq = ((soc_videosoc_uart_pending_w[0] & soc_videosoc_uart_storage[0]) | (soc_videosoc_uart_pending_w[1] & soc_videosoc_uart_storage[1]));
assign soc_videosoc_uart_tx_status = soc_videosoc_uart_tx_trigger;
assign soc_videosoc_uart_rx_status = soc_videosoc_uart_rx_trigger;
assign soc_videosoc_uart_tx_fifo_syncfifo_din = {soc_videosoc_uart_tx_fifo_fifo_in_last, soc_videosoc_uart_tx_fifo_fifo_in_first, soc_videosoc_uart_tx_fifo_fifo_in_payload_data};
assign {soc_videosoc_uart_tx_fifo_fifo_out_last, soc_videosoc_uart_tx_fifo_fifo_out_first, soc_videosoc_uart_tx_fifo_fifo_out_payload_data} = soc_videosoc_uart_tx_fifo_syncfifo_dout;
assign soc_videosoc_uart_tx_fifo_sink_ready = soc_videosoc_uart_tx_fifo_syncfifo_writable;
assign soc_videosoc_uart_tx_fifo_syncfifo_we = soc_videosoc_uart_tx_fifo_sink_valid;
assign soc_videosoc_uart_tx_fifo_fifo_in_first = soc_videosoc_uart_tx_fifo_sink_first;
assign soc_videosoc_uart_tx_fifo_fifo_in_last = soc_videosoc_uart_tx_fifo_sink_last;
assign soc_videosoc_uart_tx_fifo_fifo_in_payload_data = soc_videosoc_uart_tx_fifo_sink_payload_data;
assign soc_videosoc_uart_tx_fifo_source_valid = soc_videosoc_uart_tx_fifo_syncfifo_readable;
assign soc_videosoc_uart_tx_fifo_source_first = soc_videosoc_uart_tx_fifo_fifo_out_first;
assign soc_videosoc_uart_tx_fifo_source_last = soc_videosoc_uart_tx_fifo_fifo_out_last;
assign soc_videosoc_uart_tx_fifo_source_payload_data = soc_videosoc_uart_tx_fifo_fifo_out_payload_data;
assign soc_videosoc_uart_tx_fifo_syncfifo_re = soc_videosoc_uart_tx_fifo_source_ready;
always @(*) begin
	soc_videosoc_uart_tx_fifo_wrport_adr <= 4'd0;
	if (soc_videosoc_uart_tx_fifo_replace) begin
		soc_videosoc_uart_tx_fifo_wrport_adr <= (soc_videosoc_uart_tx_fifo_produce - 1'd1);
	end else begin
		soc_videosoc_uart_tx_fifo_wrport_adr <= soc_videosoc_uart_tx_fifo_produce;
	end
end
assign soc_videosoc_uart_tx_fifo_wrport_dat_w = soc_videosoc_uart_tx_fifo_syncfifo_din;
assign soc_videosoc_uart_tx_fifo_wrport_we = (soc_videosoc_uart_tx_fifo_syncfifo_we & (soc_videosoc_uart_tx_fifo_syncfifo_writable | soc_videosoc_uart_tx_fifo_replace));
assign soc_videosoc_uart_tx_fifo_do_read = (soc_videosoc_uart_tx_fifo_syncfifo_readable & soc_videosoc_uart_tx_fifo_syncfifo_re);
assign soc_videosoc_uart_tx_fifo_rdport_adr = soc_videosoc_uart_tx_fifo_consume;
assign soc_videosoc_uart_tx_fifo_syncfifo_dout = soc_videosoc_uart_tx_fifo_rdport_dat_r;
assign soc_videosoc_uart_tx_fifo_syncfifo_writable = (soc_videosoc_uart_tx_fifo_level != 5'd16);
assign soc_videosoc_uart_tx_fifo_syncfifo_readable = (soc_videosoc_uart_tx_fifo_level != 1'd0);
assign soc_videosoc_uart_rx_fifo_syncfifo_din = {soc_videosoc_uart_rx_fifo_fifo_in_last, soc_videosoc_uart_rx_fifo_fifo_in_first, soc_videosoc_uart_rx_fifo_fifo_in_payload_data};
assign {soc_videosoc_uart_rx_fifo_fifo_out_last, soc_videosoc_uart_rx_fifo_fifo_out_first, soc_videosoc_uart_rx_fifo_fifo_out_payload_data} = soc_videosoc_uart_rx_fifo_syncfifo_dout;
assign soc_videosoc_uart_rx_fifo_sink_ready = soc_videosoc_uart_rx_fifo_syncfifo_writable;
assign soc_videosoc_uart_rx_fifo_syncfifo_we = soc_videosoc_uart_rx_fifo_sink_valid;
assign soc_videosoc_uart_rx_fifo_fifo_in_first = soc_videosoc_uart_rx_fifo_sink_first;
assign soc_videosoc_uart_rx_fifo_fifo_in_last = soc_videosoc_uart_rx_fifo_sink_last;
assign soc_videosoc_uart_rx_fifo_fifo_in_payload_data = soc_videosoc_uart_rx_fifo_sink_payload_data;
assign soc_videosoc_uart_rx_fifo_source_valid = soc_videosoc_uart_rx_fifo_syncfifo_readable;
assign soc_videosoc_uart_rx_fifo_source_first = soc_videosoc_uart_rx_fifo_fifo_out_first;
assign soc_videosoc_uart_rx_fifo_source_last = soc_videosoc_uart_rx_fifo_fifo_out_last;
assign soc_videosoc_uart_rx_fifo_source_payload_data = soc_videosoc_uart_rx_fifo_fifo_out_payload_data;
assign soc_videosoc_uart_rx_fifo_syncfifo_re = soc_videosoc_uart_rx_fifo_source_ready;
always @(*) begin
	soc_videosoc_uart_rx_fifo_wrport_adr <= 4'd0;
	if (soc_videosoc_uart_rx_fifo_replace) begin
		soc_videosoc_uart_rx_fifo_wrport_adr <= (soc_videosoc_uart_rx_fifo_produce - 1'd1);
	end else begin
		soc_videosoc_uart_rx_fifo_wrport_adr <= soc_videosoc_uart_rx_fifo_produce;
	end
end
assign soc_videosoc_uart_rx_fifo_wrport_dat_w = soc_videosoc_uart_rx_fifo_syncfifo_din;
assign soc_videosoc_uart_rx_fifo_wrport_we = (soc_videosoc_uart_rx_fifo_syncfifo_we & (soc_videosoc_uart_rx_fifo_syncfifo_writable | soc_videosoc_uart_rx_fifo_replace));
assign soc_videosoc_uart_rx_fifo_do_read = (soc_videosoc_uart_rx_fifo_syncfifo_readable & soc_videosoc_uart_rx_fifo_syncfifo_re);
assign soc_videosoc_uart_rx_fifo_rdport_adr = soc_videosoc_uart_rx_fifo_consume;
assign soc_videosoc_uart_rx_fifo_syncfifo_dout = soc_videosoc_uart_rx_fifo_rdport_dat_r;
assign soc_videosoc_uart_rx_fifo_syncfifo_writable = (soc_videosoc_uart_rx_fifo_level != 5'd16);
assign soc_videosoc_uart_rx_fifo_syncfifo_readable = (soc_videosoc_uart_rx_fifo_level != 1'd0);
assign soc_videosoc_bridge_reset = soc_videosoc_bridge_done;
assign soc_videosoc_rs232phyinterface1_source_ready = 1'd1;
assign soc_videosoc_bridge_wishbone_adr = (soc_videosoc_bridge_address + soc_videosoc_bridge_word_counter);
assign soc_videosoc_bridge_wishbone_dat_w = soc_videosoc_bridge_data;
assign soc_videosoc_bridge_wishbone_sel = 4'd15;
always @(*) begin
	soc_videosoc_rs232phyinterface1_sink_payload_data <= 8'd0;
	case (soc_videosoc_bridge_byte_counter)
		1'd0: begin
			soc_videosoc_rs232phyinterface1_sink_payload_data <= soc_videosoc_bridge_data[31:24];
		end
		1'd1: begin
			soc_videosoc_rs232phyinterface1_sink_payload_data <= soc_videosoc_bridge_data[23:16];
		end
		2'd2: begin
			soc_videosoc_rs232phyinterface1_sink_payload_data <= soc_videosoc_bridge_data[15:8];
		end
		default: begin
			soc_videosoc_rs232phyinterface1_sink_payload_data <= soc_videosoc_bridge_data[7:0];
		end
	endcase
end
assign soc_videosoc_bridge_wait = (~soc_videosoc_bridge_is_ongoing);
assign soc_videosoc_rs232phyinterface1_sink_last = ((soc_videosoc_bridge_byte_counter == 2'd3) & (soc_videosoc_bridge_word_counter == (soc_videosoc_bridge_length - 1'd1)));
always @(*) begin
	soc_videosoc_bridge_is_ongoing <= 1'd0;
	soc_videosoc_bridge_wishbone_cyc <= 1'd0;
	soc_videosoc_bridge_wishbone_stb <= 1'd0;
	soc_videosoc_bridge_cmd_ce <= 1'd0;
	soc_videosoc_bridge_length_ce <= 1'd0;
	soc_videosoc_bridge_wishbone_we <= 1'd0;
	soc_videosoc_bridge_address_ce <= 1'd0;
	soc_videosoc_rs232phyinterface1_sink_valid <= 1'd0;
	soc_videosoc_bridge_rx_data_ce <= 1'd0;
	soc_videosoc_bridge_byte_counter_reset <= 1'd0;
	soc_videosoc_bridge_tx_data_ce <= 1'd0;
	soc_videosoc_bridge_byte_counter_ce <= 1'd0;
	vns_wishbonestreamingbridge_next_state <= 3'd0;
	soc_videosoc_bridge_word_counter_reset <= 1'd0;
	soc_videosoc_bridge_word_counter_ce <= 1'd0;
	vns_wishbonestreamingbridge_next_state <= vns_wishbonestreamingbridge_state;
	case (vns_wishbonestreamingbridge_state)
		1'd1: begin
			if (soc_videosoc_rs232phyinterface1_source_valid) begin
				soc_videosoc_bridge_length_ce <= 1'd1;
				vns_wishbonestreamingbridge_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if (soc_videosoc_rs232phyinterface1_source_valid) begin
				soc_videosoc_bridge_address_ce <= 1'd1;
				soc_videosoc_bridge_byte_counter_ce <= 1'd1;
				if ((soc_videosoc_bridge_byte_counter == 2'd3)) begin
					if ((soc_videosoc_bridge_cmd == 1'd1)) begin
						vns_wishbonestreamingbridge_next_state <= 2'd3;
					end else begin
						if ((soc_videosoc_bridge_cmd == 2'd2)) begin
							vns_wishbonestreamingbridge_next_state <= 3'd5;
						end
					end
					soc_videosoc_bridge_byte_counter_reset <= 1'd1;
				end
			end
		end
		2'd3: begin
			if (soc_videosoc_rs232phyinterface1_source_valid) begin
				soc_videosoc_bridge_rx_data_ce <= 1'd1;
				soc_videosoc_bridge_byte_counter_ce <= 1'd1;
				if ((soc_videosoc_bridge_byte_counter == 2'd3)) begin
					vns_wishbonestreamingbridge_next_state <= 3'd4;
					soc_videosoc_bridge_byte_counter_reset <= 1'd1;
				end
			end
		end
		3'd4: begin
			soc_videosoc_bridge_wishbone_stb <= 1'd1;
			soc_videosoc_bridge_wishbone_we <= 1'd1;
			soc_videosoc_bridge_wishbone_cyc <= 1'd1;
			if (soc_videosoc_bridge_wishbone_ack) begin
				soc_videosoc_bridge_word_counter_ce <= 1'd1;
				if ((soc_videosoc_bridge_word_counter == (soc_videosoc_bridge_length - 1'd1))) begin
					vns_wishbonestreamingbridge_next_state <= 1'd0;
				end else begin
					vns_wishbonestreamingbridge_next_state <= 2'd3;
				end
			end
		end
		3'd5: begin
			soc_videosoc_bridge_wishbone_stb <= 1'd1;
			soc_videosoc_bridge_wishbone_we <= 1'd0;
			soc_videosoc_bridge_wishbone_cyc <= 1'd1;
			if (soc_videosoc_bridge_wishbone_ack) begin
				soc_videosoc_bridge_tx_data_ce <= 1'd1;
				vns_wishbonestreamingbridge_next_state <= 3'd6;
			end
		end
		3'd6: begin
			soc_videosoc_rs232phyinterface1_sink_valid <= 1'd1;
			if (soc_videosoc_rs232phyinterface1_sink_ready) begin
				soc_videosoc_bridge_byte_counter_ce <= 1'd1;
				if ((soc_videosoc_bridge_byte_counter == 2'd3)) begin
					soc_videosoc_bridge_word_counter_ce <= 1'd1;
					if ((soc_videosoc_bridge_word_counter == (soc_videosoc_bridge_length - 1'd1))) begin
						vns_wishbonestreamingbridge_next_state <= 1'd0;
					end else begin
						vns_wishbonestreamingbridge_next_state <= 3'd5;
						soc_videosoc_bridge_byte_counter_reset <= 1'd1;
					end
				end
			end
		end
		default: begin
			if (soc_videosoc_rs232phyinterface1_source_valid) begin
				soc_videosoc_bridge_cmd_ce <= 1'd1;
				if (((soc_videosoc_rs232phyinterface1_source_payload_data == 1'd1) | (soc_videosoc_rs232phyinterface1_source_payload_data == 2'd2))) begin
					vns_wishbonestreamingbridge_next_state <= 1'd1;
				end
				soc_videosoc_bridge_byte_counter_reset <= 1'd1;
				soc_videosoc_bridge_word_counter_reset <= 1'd1;
			end
			soc_videosoc_bridge_is_ongoing <= 1'd1;
		end
	endcase
end
assign soc_videosoc_bridge_done = (soc_videosoc_bridge_count == 1'd0);
always @(*) begin
	soc_videosoc_rs232phyinterface0_source_valid <= 1'd0;
	soc_videosoc_uart_phy_source_ready <= 1'd0;
	soc_videosoc_rs232phyinterface0_source_first <= 1'd0;
	soc_videosoc_rs232phyinterface0_source_last <= 1'd0;
	soc_videosoc_rs232phyinterface0_source_payload_data <= 8'd0;
	soc_videosoc_rs232phyinterface1_sink_ready <= 1'd0;
	soc_videosoc_rs232phyinterface1_source_first <= 1'd0;
	soc_videosoc_uart_phy_sink_valid <= 1'd0;
	soc_videosoc_uart_phy_sink_first <= 1'd0;
	soc_videosoc_rs232phyinterface1_source_valid <= 1'd0;
	soc_videosoc_uart_phy_sink_last <= 1'd0;
	soc_videosoc_uart_phy_sink_payload_data <= 8'd0;
	soc_videosoc_rs232phyinterface0_sink_ready <= 1'd0;
	soc_videosoc_rs232phyinterface1_source_last <= 1'd0;
	soc_videosoc_rs232phyinterface1_source_payload_data <= 8'd0;
	soc_videosoc_rs232phyinterface0_sink_ready <= 1'd1;
	soc_videosoc_rs232phyinterface1_sink_ready <= 1'd1;
	case (soc_videosoc_sel)
		1'd0: begin
			soc_videosoc_rs232phyinterface0_source_valid <= soc_videosoc_uart_phy_source_valid;
			soc_videosoc_uart_phy_source_ready <= soc_videosoc_rs232phyinterface0_source_ready;
			soc_videosoc_rs232phyinterface0_source_first <= soc_videosoc_uart_phy_source_first;
			soc_videosoc_rs232phyinterface0_source_last <= soc_videosoc_uart_phy_source_last;
			soc_videosoc_rs232phyinterface0_source_payload_data <= soc_videosoc_uart_phy_source_payload_data;
			soc_videosoc_uart_phy_sink_valid <= soc_videosoc_rs232phyinterface0_sink_valid;
			soc_videosoc_rs232phyinterface0_sink_ready <= soc_videosoc_uart_phy_sink_ready;
			soc_videosoc_uart_phy_sink_first <= soc_videosoc_rs232phyinterface0_sink_first;
			soc_videosoc_uart_phy_sink_last <= soc_videosoc_rs232phyinterface0_sink_last;
			soc_videosoc_uart_phy_sink_payload_data <= soc_videosoc_rs232phyinterface0_sink_payload_data;
		end
		1'd1: begin
			soc_videosoc_rs232phyinterface1_source_valid <= soc_videosoc_uart_phy_source_valid;
			soc_videosoc_uart_phy_source_ready <= soc_videosoc_rs232phyinterface1_source_ready;
			soc_videosoc_rs232phyinterface1_source_first <= soc_videosoc_uart_phy_source_first;
			soc_videosoc_rs232phyinterface1_source_last <= soc_videosoc_uart_phy_source_last;
			soc_videosoc_rs232phyinterface1_source_payload_data <= soc_videosoc_uart_phy_source_payload_data;
			soc_videosoc_uart_phy_sink_valid <= soc_videosoc_rs232phyinterface1_sink_valid;
			soc_videosoc_rs232phyinterface1_sink_ready <= soc_videosoc_uart_phy_sink_ready;
			soc_videosoc_uart_phy_sink_first <= soc_videosoc_rs232phyinterface1_sink_first;
			soc_videosoc_uart_phy_sink_last <= soc_videosoc_rs232phyinterface1_sink_last;
			soc_videosoc_uart_phy_sink_payload_data <= soc_videosoc_rs232phyinterface1_sink_payload_data;
		end
	endcase
end
assign soc_videosoc_info_git_status = 160'd924460433538070016718210670148164609158715308002;
assign soc_videosoc_info_platform_status = 63'd7954896779841861225;
assign soc_videosoc_info_target_status = 63'd8532461355846860800;
assign oled_sclk = soc_videosoc_oled_spi_pads_clk;
assign oled_sdin = soc_videosoc_oled_spi_pads_mosi;
assign soc_videosoc_oled_spimaster_start = (soc_videosoc_oled_spimaster_ctrl_re & soc_videosoc_oled_spimaster_ctrl_r);
assign soc_videosoc_oled_spimaster_status = soc_videosoc_oled_spimaster_done;
assign soc_videosoc_oled_spimaster_set_clk = (soc_videosoc_oled_spimaster_i == 3'd7);
assign soc_videosoc_oled_spimaster_clr_clk = (soc_videosoc_oled_spimaster_i == 4'd15);
assign soc_videosoc_oled_spi_pads_cs_n = (~soc_videosoc_oled_spimaster_enable_cs);
always @(*) begin
	soc_videosoc_oled_spimaster_enable_shift <= 1'd0;
	vns_oled_next_state <= 2'd0;
	soc_videosoc_oled_spimaster_done <= 1'd0;
	soc_videosoc_oled_spimaster_clr_cnt <= 1'd0;
	soc_videosoc_oled_spimaster_inc_cnt <= 1'd0;
	soc_videosoc_oled_spimaster_irq <= 1'd0;
	soc_videosoc_oled_spimaster_enable_cs <= 1'd0;
	vns_oled_next_state <= vns_oled_state;
	case (vns_oled_state)
		1'd1: begin
			if (soc_videosoc_oled_spimaster_clr_clk) begin
				vns_oled_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if ((soc_videosoc_oled_spimaster_cnt == soc_videosoc_oled_spimaster_length_storage)) begin
				vns_oled_next_state <= 2'd3;
			end else begin
				soc_videosoc_oled_spimaster_inc_cnt <= soc_videosoc_oled_spimaster_clr_clk;
			end
			soc_videosoc_oled_spimaster_enable_cs <= 1'd1;
			soc_videosoc_oled_spimaster_enable_shift <= 1'd1;
		end
		2'd3: begin
			if (soc_videosoc_oled_spimaster_set_clk) begin
				vns_oled_next_state <= 1'd0;
			end
			soc_videosoc_oled_spimaster_enable_shift <= 1'd1;
			soc_videosoc_oled_spimaster_irq <= 1'd1;
		end
		default: begin
			if (soc_videosoc_oled_spimaster_start) begin
				vns_oled_next_state <= 1'd1;
			end
			soc_videosoc_oled_spimaster_done <= 1'd1;
			soc_videosoc_oled_spimaster_clr_cnt <= 1'd1;
		end
	endcase
end
assign {oled_vdd, oled_vbat, oled_dc, oled_res} = soc_videosoc_oled_storage;
assign soc_videosoc_ddrphy_oe = ((soc_videosoc_ddrphy_last_wrdata_en[1] | soc_videosoc_ddrphy_last_wrdata_en[2]) | soc_videosoc_ddrphy_last_wrdata_en[3]);
assign soc_videosoc_ddrphy_dfi_p0_address = soc_videosoc_sdram_master_p0_address;
assign soc_videosoc_ddrphy_dfi_p0_bank = soc_videosoc_sdram_master_p0_bank;
assign soc_videosoc_ddrphy_dfi_p0_cas_n = soc_videosoc_sdram_master_p0_cas_n;
assign soc_videosoc_ddrphy_dfi_p0_cs_n = soc_videosoc_sdram_master_p0_cs_n;
assign soc_videosoc_ddrphy_dfi_p0_ras_n = soc_videosoc_sdram_master_p0_ras_n;
assign soc_videosoc_ddrphy_dfi_p0_we_n = soc_videosoc_sdram_master_p0_we_n;
assign soc_videosoc_ddrphy_dfi_p0_cke = soc_videosoc_sdram_master_p0_cke;
assign soc_videosoc_ddrphy_dfi_p0_odt = soc_videosoc_sdram_master_p0_odt;
assign soc_videosoc_ddrphy_dfi_p0_reset_n = soc_videosoc_sdram_master_p0_reset_n;
assign soc_videosoc_ddrphy_dfi_p0_wrdata = soc_videosoc_sdram_master_p0_wrdata;
assign soc_videosoc_ddrphy_dfi_p0_wrdata_en = soc_videosoc_sdram_master_p0_wrdata_en;
assign soc_videosoc_ddrphy_dfi_p0_wrdata_mask = soc_videosoc_sdram_master_p0_wrdata_mask;
assign soc_videosoc_ddrphy_dfi_p0_rddata_en = soc_videosoc_sdram_master_p0_rddata_en;
assign soc_videosoc_sdram_master_p0_rddata = soc_videosoc_ddrphy_dfi_p0_rddata;
assign soc_videosoc_sdram_master_p0_rddata_valid = soc_videosoc_ddrphy_dfi_p0_rddata_valid;
assign soc_videosoc_ddrphy_dfi_p1_address = soc_videosoc_sdram_master_p1_address;
assign soc_videosoc_ddrphy_dfi_p1_bank = soc_videosoc_sdram_master_p1_bank;
assign soc_videosoc_ddrphy_dfi_p1_cas_n = soc_videosoc_sdram_master_p1_cas_n;
assign soc_videosoc_ddrphy_dfi_p1_cs_n = soc_videosoc_sdram_master_p1_cs_n;
assign soc_videosoc_ddrphy_dfi_p1_ras_n = soc_videosoc_sdram_master_p1_ras_n;
assign soc_videosoc_ddrphy_dfi_p1_we_n = soc_videosoc_sdram_master_p1_we_n;
assign soc_videosoc_ddrphy_dfi_p1_cke = soc_videosoc_sdram_master_p1_cke;
assign soc_videosoc_ddrphy_dfi_p1_odt = soc_videosoc_sdram_master_p1_odt;
assign soc_videosoc_ddrphy_dfi_p1_reset_n = soc_videosoc_sdram_master_p1_reset_n;
assign soc_videosoc_ddrphy_dfi_p1_wrdata = soc_videosoc_sdram_master_p1_wrdata;
assign soc_videosoc_ddrphy_dfi_p1_wrdata_en = soc_videosoc_sdram_master_p1_wrdata_en;
assign soc_videosoc_ddrphy_dfi_p1_wrdata_mask = soc_videosoc_sdram_master_p1_wrdata_mask;
assign soc_videosoc_ddrphy_dfi_p1_rddata_en = soc_videosoc_sdram_master_p1_rddata_en;
assign soc_videosoc_sdram_master_p1_rddata = soc_videosoc_ddrphy_dfi_p1_rddata;
assign soc_videosoc_sdram_master_p1_rddata_valid = soc_videosoc_ddrphy_dfi_p1_rddata_valid;
assign soc_videosoc_ddrphy_dfi_p2_address = soc_videosoc_sdram_master_p2_address;
assign soc_videosoc_ddrphy_dfi_p2_bank = soc_videosoc_sdram_master_p2_bank;
assign soc_videosoc_ddrphy_dfi_p2_cas_n = soc_videosoc_sdram_master_p2_cas_n;
assign soc_videosoc_ddrphy_dfi_p2_cs_n = soc_videosoc_sdram_master_p2_cs_n;
assign soc_videosoc_ddrphy_dfi_p2_ras_n = soc_videosoc_sdram_master_p2_ras_n;
assign soc_videosoc_ddrphy_dfi_p2_we_n = soc_videosoc_sdram_master_p2_we_n;
assign soc_videosoc_ddrphy_dfi_p2_cke = soc_videosoc_sdram_master_p2_cke;
assign soc_videosoc_ddrphy_dfi_p2_odt = soc_videosoc_sdram_master_p2_odt;
assign soc_videosoc_ddrphy_dfi_p2_reset_n = soc_videosoc_sdram_master_p2_reset_n;
assign soc_videosoc_ddrphy_dfi_p2_wrdata = soc_videosoc_sdram_master_p2_wrdata;
assign soc_videosoc_ddrphy_dfi_p2_wrdata_en = soc_videosoc_sdram_master_p2_wrdata_en;
assign soc_videosoc_ddrphy_dfi_p2_wrdata_mask = soc_videosoc_sdram_master_p2_wrdata_mask;
assign soc_videosoc_ddrphy_dfi_p2_rddata_en = soc_videosoc_sdram_master_p2_rddata_en;
assign soc_videosoc_sdram_master_p2_rddata = soc_videosoc_ddrphy_dfi_p2_rddata;
assign soc_videosoc_sdram_master_p2_rddata_valid = soc_videosoc_ddrphy_dfi_p2_rddata_valid;
assign soc_videosoc_ddrphy_dfi_p3_address = soc_videosoc_sdram_master_p3_address;
assign soc_videosoc_ddrphy_dfi_p3_bank = soc_videosoc_sdram_master_p3_bank;
assign soc_videosoc_ddrphy_dfi_p3_cas_n = soc_videosoc_sdram_master_p3_cas_n;
assign soc_videosoc_ddrphy_dfi_p3_cs_n = soc_videosoc_sdram_master_p3_cs_n;
assign soc_videosoc_ddrphy_dfi_p3_ras_n = soc_videosoc_sdram_master_p3_ras_n;
assign soc_videosoc_ddrphy_dfi_p3_we_n = soc_videosoc_sdram_master_p3_we_n;
assign soc_videosoc_ddrphy_dfi_p3_cke = soc_videosoc_sdram_master_p3_cke;
assign soc_videosoc_ddrphy_dfi_p3_odt = soc_videosoc_sdram_master_p3_odt;
assign soc_videosoc_ddrphy_dfi_p3_reset_n = soc_videosoc_sdram_master_p3_reset_n;
assign soc_videosoc_ddrphy_dfi_p3_wrdata = soc_videosoc_sdram_master_p3_wrdata;
assign soc_videosoc_ddrphy_dfi_p3_wrdata_en = soc_videosoc_sdram_master_p3_wrdata_en;
assign soc_videosoc_ddrphy_dfi_p3_wrdata_mask = soc_videosoc_sdram_master_p3_wrdata_mask;
assign soc_videosoc_ddrphy_dfi_p3_rddata_en = soc_videosoc_sdram_master_p3_rddata_en;
assign soc_videosoc_sdram_master_p3_rddata = soc_videosoc_ddrphy_dfi_p3_rddata;
assign soc_videosoc_sdram_master_p3_rddata_valid = soc_videosoc_ddrphy_dfi_p3_rddata_valid;
assign soc_videosoc_sdram_slave_p0_address = soc_videosoc_sdram_dfi_p0_address;
assign soc_videosoc_sdram_slave_p0_bank = soc_videosoc_sdram_dfi_p0_bank;
assign soc_videosoc_sdram_slave_p0_cas_n = soc_videosoc_sdram_dfi_p0_cas_n;
assign soc_videosoc_sdram_slave_p0_cs_n = soc_videosoc_sdram_dfi_p0_cs_n;
assign soc_videosoc_sdram_slave_p0_ras_n = soc_videosoc_sdram_dfi_p0_ras_n;
assign soc_videosoc_sdram_slave_p0_we_n = soc_videosoc_sdram_dfi_p0_we_n;
assign soc_videosoc_sdram_slave_p0_cke = soc_videosoc_sdram_dfi_p0_cke;
assign soc_videosoc_sdram_slave_p0_odt = soc_videosoc_sdram_dfi_p0_odt;
assign soc_videosoc_sdram_slave_p0_reset_n = soc_videosoc_sdram_dfi_p0_reset_n;
assign soc_videosoc_sdram_slave_p0_wrdata = soc_videosoc_sdram_dfi_p0_wrdata;
assign soc_videosoc_sdram_slave_p0_wrdata_en = soc_videosoc_sdram_dfi_p0_wrdata_en;
assign soc_videosoc_sdram_slave_p0_wrdata_mask = soc_videosoc_sdram_dfi_p0_wrdata_mask;
assign soc_videosoc_sdram_slave_p0_rddata_en = soc_videosoc_sdram_dfi_p0_rddata_en;
assign soc_videosoc_sdram_dfi_p0_rddata = soc_videosoc_sdram_slave_p0_rddata;
assign soc_videosoc_sdram_dfi_p0_rddata_valid = soc_videosoc_sdram_slave_p0_rddata_valid;
assign soc_videosoc_sdram_slave_p1_address = soc_videosoc_sdram_dfi_p1_address;
assign soc_videosoc_sdram_slave_p1_bank = soc_videosoc_sdram_dfi_p1_bank;
assign soc_videosoc_sdram_slave_p1_cas_n = soc_videosoc_sdram_dfi_p1_cas_n;
assign soc_videosoc_sdram_slave_p1_cs_n = soc_videosoc_sdram_dfi_p1_cs_n;
assign soc_videosoc_sdram_slave_p1_ras_n = soc_videosoc_sdram_dfi_p1_ras_n;
assign soc_videosoc_sdram_slave_p1_we_n = soc_videosoc_sdram_dfi_p1_we_n;
assign soc_videosoc_sdram_slave_p1_cke = soc_videosoc_sdram_dfi_p1_cke;
assign soc_videosoc_sdram_slave_p1_odt = soc_videosoc_sdram_dfi_p1_odt;
assign soc_videosoc_sdram_slave_p1_reset_n = soc_videosoc_sdram_dfi_p1_reset_n;
assign soc_videosoc_sdram_slave_p1_wrdata = soc_videosoc_sdram_dfi_p1_wrdata;
assign soc_videosoc_sdram_slave_p1_wrdata_en = soc_videosoc_sdram_dfi_p1_wrdata_en;
assign soc_videosoc_sdram_slave_p1_wrdata_mask = soc_videosoc_sdram_dfi_p1_wrdata_mask;
assign soc_videosoc_sdram_slave_p1_rddata_en = soc_videosoc_sdram_dfi_p1_rddata_en;
assign soc_videosoc_sdram_dfi_p1_rddata = soc_videosoc_sdram_slave_p1_rddata;
assign soc_videosoc_sdram_dfi_p1_rddata_valid = soc_videosoc_sdram_slave_p1_rddata_valid;
assign soc_videosoc_sdram_slave_p2_address = soc_videosoc_sdram_dfi_p2_address;
assign soc_videosoc_sdram_slave_p2_bank = soc_videosoc_sdram_dfi_p2_bank;
assign soc_videosoc_sdram_slave_p2_cas_n = soc_videosoc_sdram_dfi_p2_cas_n;
assign soc_videosoc_sdram_slave_p2_cs_n = soc_videosoc_sdram_dfi_p2_cs_n;
assign soc_videosoc_sdram_slave_p2_ras_n = soc_videosoc_sdram_dfi_p2_ras_n;
assign soc_videosoc_sdram_slave_p2_we_n = soc_videosoc_sdram_dfi_p2_we_n;
assign soc_videosoc_sdram_slave_p2_cke = soc_videosoc_sdram_dfi_p2_cke;
assign soc_videosoc_sdram_slave_p2_odt = soc_videosoc_sdram_dfi_p2_odt;
assign soc_videosoc_sdram_slave_p2_reset_n = soc_videosoc_sdram_dfi_p2_reset_n;
assign soc_videosoc_sdram_slave_p2_wrdata = soc_videosoc_sdram_dfi_p2_wrdata;
assign soc_videosoc_sdram_slave_p2_wrdata_en = soc_videosoc_sdram_dfi_p2_wrdata_en;
assign soc_videosoc_sdram_slave_p2_wrdata_mask = soc_videosoc_sdram_dfi_p2_wrdata_mask;
assign soc_videosoc_sdram_slave_p2_rddata_en = soc_videosoc_sdram_dfi_p2_rddata_en;
assign soc_videosoc_sdram_dfi_p2_rddata = soc_videosoc_sdram_slave_p2_rddata;
assign soc_videosoc_sdram_dfi_p2_rddata_valid = soc_videosoc_sdram_slave_p2_rddata_valid;
assign soc_videosoc_sdram_slave_p3_address = soc_videosoc_sdram_dfi_p3_address;
assign soc_videosoc_sdram_slave_p3_bank = soc_videosoc_sdram_dfi_p3_bank;
assign soc_videosoc_sdram_slave_p3_cas_n = soc_videosoc_sdram_dfi_p3_cas_n;
assign soc_videosoc_sdram_slave_p3_cs_n = soc_videosoc_sdram_dfi_p3_cs_n;
assign soc_videosoc_sdram_slave_p3_ras_n = soc_videosoc_sdram_dfi_p3_ras_n;
assign soc_videosoc_sdram_slave_p3_we_n = soc_videosoc_sdram_dfi_p3_we_n;
assign soc_videosoc_sdram_slave_p3_cke = soc_videosoc_sdram_dfi_p3_cke;
assign soc_videosoc_sdram_slave_p3_odt = soc_videosoc_sdram_dfi_p3_odt;
assign soc_videosoc_sdram_slave_p3_reset_n = soc_videosoc_sdram_dfi_p3_reset_n;
assign soc_videosoc_sdram_slave_p3_wrdata = soc_videosoc_sdram_dfi_p3_wrdata;
assign soc_videosoc_sdram_slave_p3_wrdata_en = soc_videosoc_sdram_dfi_p3_wrdata_en;
assign soc_videosoc_sdram_slave_p3_wrdata_mask = soc_videosoc_sdram_dfi_p3_wrdata_mask;
assign soc_videosoc_sdram_slave_p3_rddata_en = soc_videosoc_sdram_dfi_p3_rddata_en;
assign soc_videosoc_sdram_dfi_p3_rddata = soc_videosoc_sdram_slave_p3_rddata;
assign soc_videosoc_sdram_dfi_p3_rddata_valid = soc_videosoc_sdram_slave_p3_rddata_valid;
always @(*) begin
	soc_videosoc_sdram_master_p2_cs_n <= 1'd1;
	soc_videosoc_sdram_master_p2_ras_n <= 1'd1;
	soc_videosoc_sdram_master_p2_we_n <= 1'd1;
	soc_videosoc_sdram_inti_p2_rddata <= 32'd0;
	soc_videosoc_sdram_master_p2_cke <= 1'd0;
	soc_videosoc_sdram_inti_p2_rddata_valid <= 1'd0;
	soc_videosoc_sdram_master_p2_odt <= 1'd0;
	soc_videosoc_sdram_master_p2_reset_n <= 1'd0;
	soc_videosoc_sdram_master_p2_wrdata <= 32'd0;
	soc_videosoc_sdram_master_p2_wrdata_en <= 1'd0;
	soc_videosoc_sdram_master_p2_wrdata_mask <= 4'd0;
	soc_videosoc_sdram_master_p2_rddata_en <= 1'd0;
	soc_videosoc_sdram_master_p3_address <= 15'd0;
	soc_videosoc_sdram_master_p3_bank <= 3'd0;
	soc_videosoc_sdram_master_p3_cas_n <= 1'd1;
	soc_videosoc_sdram_master_p3_cs_n <= 1'd1;
	soc_videosoc_sdram_master_p3_ras_n <= 1'd1;
	soc_videosoc_sdram_master_p3_we_n <= 1'd1;
	soc_videosoc_sdram_inti_p3_rddata <= 32'd0;
	soc_videosoc_sdram_master_p3_cke <= 1'd0;
	soc_videosoc_sdram_inti_p3_rddata_valid <= 1'd0;
	soc_videosoc_sdram_master_p3_odt <= 1'd0;
	soc_videosoc_sdram_master_p3_reset_n <= 1'd0;
	soc_videosoc_sdram_master_p3_wrdata <= 32'd0;
	soc_videosoc_sdram_master_p3_wrdata_en <= 1'd0;
	soc_videosoc_sdram_master_p3_wrdata_mask <= 4'd0;
	soc_videosoc_sdram_master_p3_rddata_en <= 1'd0;
	soc_videosoc_sdram_slave_p0_rddata <= 32'd0;
	soc_videosoc_sdram_slave_p0_rddata_valid <= 1'd0;
	soc_videosoc_sdram_slave_p1_rddata <= 32'd0;
	soc_videosoc_sdram_slave_p1_rddata_valid <= 1'd0;
	soc_videosoc_sdram_slave_p2_rddata <= 32'd0;
	soc_videosoc_sdram_slave_p2_rddata_valid <= 1'd0;
	soc_videosoc_sdram_slave_p3_rddata <= 32'd0;
	soc_videosoc_sdram_slave_p3_rddata_valid <= 1'd0;
	soc_videosoc_sdram_master_p0_address <= 15'd0;
	soc_videosoc_sdram_master_p0_bank <= 3'd0;
	soc_videosoc_sdram_master_p0_cas_n <= 1'd1;
	soc_videosoc_sdram_master_p0_cs_n <= 1'd1;
	soc_videosoc_sdram_master_p0_ras_n <= 1'd1;
	soc_videosoc_sdram_master_p0_we_n <= 1'd1;
	soc_videosoc_sdram_inti_p0_rddata <= 32'd0;
	soc_videosoc_sdram_master_p0_cke <= 1'd0;
	soc_videosoc_sdram_inti_p0_rddata_valid <= 1'd0;
	soc_videosoc_sdram_master_p0_odt <= 1'd0;
	soc_videosoc_sdram_master_p0_reset_n <= 1'd0;
	soc_videosoc_sdram_master_p0_wrdata <= 32'd0;
	soc_videosoc_sdram_master_p0_wrdata_en <= 1'd0;
	soc_videosoc_sdram_master_p0_wrdata_mask <= 4'd0;
	soc_videosoc_sdram_master_p0_rddata_en <= 1'd0;
	soc_videosoc_sdram_master_p1_address <= 15'd0;
	soc_videosoc_sdram_master_p1_bank <= 3'd0;
	soc_videosoc_sdram_master_p1_cas_n <= 1'd1;
	soc_videosoc_sdram_master_p1_cs_n <= 1'd1;
	soc_videosoc_sdram_master_p1_ras_n <= 1'd1;
	soc_videosoc_sdram_master_p1_we_n <= 1'd1;
	soc_videosoc_sdram_inti_p1_rddata <= 32'd0;
	soc_videosoc_sdram_master_p1_cke <= 1'd0;
	soc_videosoc_sdram_inti_p1_rddata_valid <= 1'd0;
	soc_videosoc_sdram_master_p1_odt <= 1'd0;
	soc_videosoc_sdram_master_p1_reset_n <= 1'd0;
	soc_videosoc_sdram_master_p1_wrdata <= 32'd0;
	soc_videosoc_sdram_master_p1_wrdata_en <= 1'd0;
	soc_videosoc_sdram_master_p1_wrdata_mask <= 4'd0;
	soc_videosoc_sdram_master_p1_rddata_en <= 1'd0;
	soc_videosoc_sdram_master_p2_address <= 15'd0;
	soc_videosoc_sdram_master_p2_bank <= 3'd0;
	soc_videosoc_sdram_master_p2_cas_n <= 1'd1;
	if (soc_videosoc_sdram_storage[0]) begin
		soc_videosoc_sdram_master_p0_address <= soc_videosoc_sdram_slave_p0_address;
		soc_videosoc_sdram_master_p0_bank <= soc_videosoc_sdram_slave_p0_bank;
		soc_videosoc_sdram_master_p0_cas_n <= soc_videosoc_sdram_slave_p0_cas_n;
		soc_videosoc_sdram_master_p0_cs_n <= soc_videosoc_sdram_slave_p0_cs_n;
		soc_videosoc_sdram_master_p0_ras_n <= soc_videosoc_sdram_slave_p0_ras_n;
		soc_videosoc_sdram_master_p0_we_n <= soc_videosoc_sdram_slave_p0_we_n;
		soc_videosoc_sdram_master_p0_cke <= soc_videosoc_sdram_slave_p0_cke;
		soc_videosoc_sdram_master_p0_odt <= soc_videosoc_sdram_slave_p0_odt;
		soc_videosoc_sdram_master_p0_reset_n <= soc_videosoc_sdram_slave_p0_reset_n;
		soc_videosoc_sdram_master_p0_wrdata <= soc_videosoc_sdram_slave_p0_wrdata;
		soc_videosoc_sdram_master_p0_wrdata_en <= soc_videosoc_sdram_slave_p0_wrdata_en;
		soc_videosoc_sdram_master_p0_wrdata_mask <= soc_videosoc_sdram_slave_p0_wrdata_mask;
		soc_videosoc_sdram_master_p0_rddata_en <= soc_videosoc_sdram_slave_p0_rddata_en;
		soc_videosoc_sdram_slave_p0_rddata <= soc_videosoc_sdram_master_p0_rddata;
		soc_videosoc_sdram_slave_p0_rddata_valid <= soc_videosoc_sdram_master_p0_rddata_valid;
		soc_videosoc_sdram_master_p1_address <= soc_videosoc_sdram_slave_p1_address;
		soc_videosoc_sdram_master_p1_bank <= soc_videosoc_sdram_slave_p1_bank;
		soc_videosoc_sdram_master_p1_cas_n <= soc_videosoc_sdram_slave_p1_cas_n;
		soc_videosoc_sdram_master_p1_cs_n <= soc_videosoc_sdram_slave_p1_cs_n;
		soc_videosoc_sdram_master_p1_ras_n <= soc_videosoc_sdram_slave_p1_ras_n;
		soc_videosoc_sdram_master_p1_we_n <= soc_videosoc_sdram_slave_p1_we_n;
		soc_videosoc_sdram_master_p1_cke <= soc_videosoc_sdram_slave_p1_cke;
		soc_videosoc_sdram_master_p1_odt <= soc_videosoc_sdram_slave_p1_odt;
		soc_videosoc_sdram_master_p1_reset_n <= soc_videosoc_sdram_slave_p1_reset_n;
		soc_videosoc_sdram_master_p1_wrdata <= soc_videosoc_sdram_slave_p1_wrdata;
		soc_videosoc_sdram_master_p1_wrdata_en <= soc_videosoc_sdram_slave_p1_wrdata_en;
		soc_videosoc_sdram_master_p1_wrdata_mask <= soc_videosoc_sdram_slave_p1_wrdata_mask;
		soc_videosoc_sdram_master_p1_rddata_en <= soc_videosoc_sdram_slave_p1_rddata_en;
		soc_videosoc_sdram_slave_p1_rddata <= soc_videosoc_sdram_master_p1_rddata;
		soc_videosoc_sdram_slave_p1_rddata_valid <= soc_videosoc_sdram_master_p1_rddata_valid;
		soc_videosoc_sdram_master_p2_address <= soc_videosoc_sdram_slave_p2_address;
		soc_videosoc_sdram_master_p2_bank <= soc_videosoc_sdram_slave_p2_bank;
		soc_videosoc_sdram_master_p2_cas_n <= soc_videosoc_sdram_slave_p2_cas_n;
		soc_videosoc_sdram_master_p2_cs_n <= soc_videosoc_sdram_slave_p2_cs_n;
		soc_videosoc_sdram_master_p2_ras_n <= soc_videosoc_sdram_slave_p2_ras_n;
		soc_videosoc_sdram_master_p2_we_n <= soc_videosoc_sdram_slave_p2_we_n;
		soc_videosoc_sdram_master_p2_cke <= soc_videosoc_sdram_slave_p2_cke;
		soc_videosoc_sdram_master_p2_odt <= soc_videosoc_sdram_slave_p2_odt;
		soc_videosoc_sdram_master_p2_reset_n <= soc_videosoc_sdram_slave_p2_reset_n;
		soc_videosoc_sdram_master_p2_wrdata <= soc_videosoc_sdram_slave_p2_wrdata;
		soc_videosoc_sdram_master_p2_wrdata_en <= soc_videosoc_sdram_slave_p2_wrdata_en;
		soc_videosoc_sdram_master_p2_wrdata_mask <= soc_videosoc_sdram_slave_p2_wrdata_mask;
		soc_videosoc_sdram_master_p2_rddata_en <= soc_videosoc_sdram_slave_p2_rddata_en;
		soc_videosoc_sdram_slave_p2_rddata <= soc_videosoc_sdram_master_p2_rddata;
		soc_videosoc_sdram_slave_p2_rddata_valid <= soc_videosoc_sdram_master_p2_rddata_valid;
		soc_videosoc_sdram_master_p3_address <= soc_videosoc_sdram_slave_p3_address;
		soc_videosoc_sdram_master_p3_bank <= soc_videosoc_sdram_slave_p3_bank;
		soc_videosoc_sdram_master_p3_cas_n <= soc_videosoc_sdram_slave_p3_cas_n;
		soc_videosoc_sdram_master_p3_cs_n <= soc_videosoc_sdram_slave_p3_cs_n;
		soc_videosoc_sdram_master_p3_ras_n <= soc_videosoc_sdram_slave_p3_ras_n;
		soc_videosoc_sdram_master_p3_we_n <= soc_videosoc_sdram_slave_p3_we_n;
		soc_videosoc_sdram_master_p3_cke <= soc_videosoc_sdram_slave_p3_cke;
		soc_videosoc_sdram_master_p3_odt <= soc_videosoc_sdram_slave_p3_odt;
		soc_videosoc_sdram_master_p3_reset_n <= soc_videosoc_sdram_slave_p3_reset_n;
		soc_videosoc_sdram_master_p3_wrdata <= soc_videosoc_sdram_slave_p3_wrdata;
		soc_videosoc_sdram_master_p3_wrdata_en <= soc_videosoc_sdram_slave_p3_wrdata_en;
		soc_videosoc_sdram_master_p3_wrdata_mask <= soc_videosoc_sdram_slave_p3_wrdata_mask;
		soc_videosoc_sdram_master_p3_rddata_en <= soc_videosoc_sdram_slave_p3_rddata_en;
		soc_videosoc_sdram_slave_p3_rddata <= soc_videosoc_sdram_master_p3_rddata;
		soc_videosoc_sdram_slave_p3_rddata_valid <= soc_videosoc_sdram_master_p3_rddata_valid;
	end else begin
		soc_videosoc_sdram_master_p0_address <= soc_videosoc_sdram_inti_p0_address;
		soc_videosoc_sdram_master_p0_bank <= soc_videosoc_sdram_inti_p0_bank;
		soc_videosoc_sdram_master_p0_cas_n <= soc_videosoc_sdram_inti_p0_cas_n;
		soc_videosoc_sdram_master_p0_cs_n <= soc_videosoc_sdram_inti_p0_cs_n;
		soc_videosoc_sdram_master_p0_ras_n <= soc_videosoc_sdram_inti_p0_ras_n;
		soc_videosoc_sdram_master_p0_we_n <= soc_videosoc_sdram_inti_p0_we_n;
		soc_videosoc_sdram_master_p0_cke <= soc_videosoc_sdram_inti_p0_cke;
		soc_videosoc_sdram_master_p0_odt <= soc_videosoc_sdram_inti_p0_odt;
		soc_videosoc_sdram_master_p0_reset_n <= soc_videosoc_sdram_inti_p0_reset_n;
		soc_videosoc_sdram_master_p0_wrdata <= soc_videosoc_sdram_inti_p0_wrdata;
		soc_videosoc_sdram_master_p0_wrdata_en <= soc_videosoc_sdram_inti_p0_wrdata_en;
		soc_videosoc_sdram_master_p0_wrdata_mask <= soc_videosoc_sdram_inti_p0_wrdata_mask;
		soc_videosoc_sdram_master_p0_rddata_en <= soc_videosoc_sdram_inti_p0_rddata_en;
		soc_videosoc_sdram_inti_p0_rddata <= soc_videosoc_sdram_master_p0_rddata;
		soc_videosoc_sdram_inti_p0_rddata_valid <= soc_videosoc_sdram_master_p0_rddata_valid;
		soc_videosoc_sdram_master_p1_address <= soc_videosoc_sdram_inti_p1_address;
		soc_videosoc_sdram_master_p1_bank <= soc_videosoc_sdram_inti_p1_bank;
		soc_videosoc_sdram_master_p1_cas_n <= soc_videosoc_sdram_inti_p1_cas_n;
		soc_videosoc_sdram_master_p1_cs_n <= soc_videosoc_sdram_inti_p1_cs_n;
		soc_videosoc_sdram_master_p1_ras_n <= soc_videosoc_sdram_inti_p1_ras_n;
		soc_videosoc_sdram_master_p1_we_n <= soc_videosoc_sdram_inti_p1_we_n;
		soc_videosoc_sdram_master_p1_cke <= soc_videosoc_sdram_inti_p1_cke;
		soc_videosoc_sdram_master_p1_odt <= soc_videosoc_sdram_inti_p1_odt;
		soc_videosoc_sdram_master_p1_reset_n <= soc_videosoc_sdram_inti_p1_reset_n;
		soc_videosoc_sdram_master_p1_wrdata <= soc_videosoc_sdram_inti_p1_wrdata;
		soc_videosoc_sdram_master_p1_wrdata_en <= soc_videosoc_sdram_inti_p1_wrdata_en;
		soc_videosoc_sdram_master_p1_wrdata_mask <= soc_videosoc_sdram_inti_p1_wrdata_mask;
		soc_videosoc_sdram_master_p1_rddata_en <= soc_videosoc_sdram_inti_p1_rddata_en;
		soc_videosoc_sdram_inti_p1_rddata <= soc_videosoc_sdram_master_p1_rddata;
		soc_videosoc_sdram_inti_p1_rddata_valid <= soc_videosoc_sdram_master_p1_rddata_valid;
		soc_videosoc_sdram_master_p2_address <= soc_videosoc_sdram_inti_p2_address;
		soc_videosoc_sdram_master_p2_bank <= soc_videosoc_sdram_inti_p2_bank;
		soc_videosoc_sdram_master_p2_cas_n <= soc_videosoc_sdram_inti_p2_cas_n;
		soc_videosoc_sdram_master_p2_cs_n <= soc_videosoc_sdram_inti_p2_cs_n;
		soc_videosoc_sdram_master_p2_ras_n <= soc_videosoc_sdram_inti_p2_ras_n;
		soc_videosoc_sdram_master_p2_we_n <= soc_videosoc_sdram_inti_p2_we_n;
		soc_videosoc_sdram_master_p2_cke <= soc_videosoc_sdram_inti_p2_cke;
		soc_videosoc_sdram_master_p2_odt <= soc_videosoc_sdram_inti_p2_odt;
		soc_videosoc_sdram_master_p2_reset_n <= soc_videosoc_sdram_inti_p2_reset_n;
		soc_videosoc_sdram_master_p2_wrdata <= soc_videosoc_sdram_inti_p2_wrdata;
		soc_videosoc_sdram_master_p2_wrdata_en <= soc_videosoc_sdram_inti_p2_wrdata_en;
		soc_videosoc_sdram_master_p2_wrdata_mask <= soc_videosoc_sdram_inti_p2_wrdata_mask;
		soc_videosoc_sdram_master_p2_rddata_en <= soc_videosoc_sdram_inti_p2_rddata_en;
		soc_videosoc_sdram_inti_p2_rddata <= soc_videosoc_sdram_master_p2_rddata;
		soc_videosoc_sdram_inti_p2_rddata_valid <= soc_videosoc_sdram_master_p2_rddata_valid;
		soc_videosoc_sdram_master_p3_address <= soc_videosoc_sdram_inti_p3_address;
		soc_videosoc_sdram_master_p3_bank <= soc_videosoc_sdram_inti_p3_bank;
		soc_videosoc_sdram_master_p3_cas_n <= soc_videosoc_sdram_inti_p3_cas_n;
		soc_videosoc_sdram_master_p3_cs_n <= soc_videosoc_sdram_inti_p3_cs_n;
		soc_videosoc_sdram_master_p3_ras_n <= soc_videosoc_sdram_inti_p3_ras_n;
		soc_videosoc_sdram_master_p3_we_n <= soc_videosoc_sdram_inti_p3_we_n;
		soc_videosoc_sdram_master_p3_cke <= soc_videosoc_sdram_inti_p3_cke;
		soc_videosoc_sdram_master_p3_odt <= soc_videosoc_sdram_inti_p3_odt;
		soc_videosoc_sdram_master_p3_reset_n <= soc_videosoc_sdram_inti_p3_reset_n;
		soc_videosoc_sdram_master_p3_wrdata <= soc_videosoc_sdram_inti_p3_wrdata;
		soc_videosoc_sdram_master_p3_wrdata_en <= soc_videosoc_sdram_inti_p3_wrdata_en;
		soc_videosoc_sdram_master_p3_wrdata_mask <= soc_videosoc_sdram_inti_p3_wrdata_mask;
		soc_videosoc_sdram_master_p3_rddata_en <= soc_videosoc_sdram_inti_p3_rddata_en;
		soc_videosoc_sdram_inti_p3_rddata <= soc_videosoc_sdram_master_p3_rddata;
		soc_videosoc_sdram_inti_p3_rddata_valid <= soc_videosoc_sdram_master_p3_rddata_valid;
	end
end
assign soc_videosoc_sdram_inti_p0_cke = soc_videosoc_sdram_storage[1];
assign soc_videosoc_sdram_inti_p1_cke = soc_videosoc_sdram_storage[1];
assign soc_videosoc_sdram_inti_p2_cke = soc_videosoc_sdram_storage[1];
assign soc_videosoc_sdram_inti_p3_cke = soc_videosoc_sdram_storage[1];
assign soc_videosoc_sdram_inti_p0_odt = soc_videosoc_sdram_storage[2];
assign soc_videosoc_sdram_inti_p1_odt = soc_videosoc_sdram_storage[2];
assign soc_videosoc_sdram_inti_p2_odt = soc_videosoc_sdram_storage[2];
assign soc_videosoc_sdram_inti_p3_odt = soc_videosoc_sdram_storage[2];
assign soc_videosoc_sdram_inti_p0_reset_n = soc_videosoc_sdram_storage[3];
assign soc_videosoc_sdram_inti_p1_reset_n = soc_videosoc_sdram_storage[3];
assign soc_videosoc_sdram_inti_p2_reset_n = soc_videosoc_sdram_storage[3];
assign soc_videosoc_sdram_inti_p3_reset_n = soc_videosoc_sdram_storage[3];
always @(*) begin
	soc_videosoc_sdram_inti_p0_we_n <= 1'd1;
	soc_videosoc_sdram_inti_p0_cas_n <= 1'd1;
	soc_videosoc_sdram_inti_p0_cs_n <= 1'd1;
	soc_videosoc_sdram_inti_p0_ras_n <= 1'd1;
	if (soc_videosoc_sdram_phaseinjector0_command_issue_re) begin
		soc_videosoc_sdram_inti_p0_cs_n <= (~soc_videosoc_sdram_phaseinjector0_command_storage[0]);
		soc_videosoc_sdram_inti_p0_we_n <= (~soc_videosoc_sdram_phaseinjector0_command_storage[1]);
		soc_videosoc_sdram_inti_p0_cas_n <= (~soc_videosoc_sdram_phaseinjector0_command_storage[2]);
		soc_videosoc_sdram_inti_p0_ras_n <= (~soc_videosoc_sdram_phaseinjector0_command_storage[3]);
	end else begin
		soc_videosoc_sdram_inti_p0_cs_n <= 1'd1;
		soc_videosoc_sdram_inti_p0_we_n <= 1'd1;
		soc_videosoc_sdram_inti_p0_cas_n <= 1'd1;
		soc_videosoc_sdram_inti_p0_ras_n <= 1'd1;
	end
end
assign soc_videosoc_sdram_inti_p0_address = soc_videosoc_sdram_phaseinjector0_address_storage;
assign soc_videosoc_sdram_inti_p0_bank = soc_videosoc_sdram_phaseinjector0_baddress_storage;
assign soc_videosoc_sdram_inti_p0_wrdata_en = (soc_videosoc_sdram_phaseinjector0_command_issue_re & soc_videosoc_sdram_phaseinjector0_command_storage[4]);
assign soc_videosoc_sdram_inti_p0_rddata_en = (soc_videosoc_sdram_phaseinjector0_command_issue_re & soc_videosoc_sdram_phaseinjector0_command_storage[5]);
assign soc_videosoc_sdram_inti_p0_wrdata = soc_videosoc_sdram_phaseinjector0_wrdata_storage;
assign soc_videosoc_sdram_inti_p0_wrdata_mask = 1'd0;
always @(*) begin
	soc_videosoc_sdram_inti_p1_cas_n <= 1'd1;
	soc_videosoc_sdram_inti_p1_cs_n <= 1'd1;
	soc_videosoc_sdram_inti_p1_ras_n <= 1'd1;
	soc_videosoc_sdram_inti_p1_we_n <= 1'd1;
	if (soc_videosoc_sdram_phaseinjector1_command_issue_re) begin
		soc_videosoc_sdram_inti_p1_cs_n <= (~soc_videosoc_sdram_phaseinjector1_command_storage[0]);
		soc_videosoc_sdram_inti_p1_we_n <= (~soc_videosoc_sdram_phaseinjector1_command_storage[1]);
		soc_videosoc_sdram_inti_p1_cas_n <= (~soc_videosoc_sdram_phaseinjector1_command_storage[2]);
		soc_videosoc_sdram_inti_p1_ras_n <= (~soc_videosoc_sdram_phaseinjector1_command_storage[3]);
	end else begin
		soc_videosoc_sdram_inti_p1_cs_n <= 1'd1;
		soc_videosoc_sdram_inti_p1_we_n <= 1'd1;
		soc_videosoc_sdram_inti_p1_cas_n <= 1'd1;
		soc_videosoc_sdram_inti_p1_ras_n <= 1'd1;
	end
end
assign soc_videosoc_sdram_inti_p1_address = soc_videosoc_sdram_phaseinjector1_address_storage;
assign soc_videosoc_sdram_inti_p1_bank = soc_videosoc_sdram_phaseinjector1_baddress_storage;
assign soc_videosoc_sdram_inti_p1_wrdata_en = (soc_videosoc_sdram_phaseinjector1_command_issue_re & soc_videosoc_sdram_phaseinjector1_command_storage[4]);
assign soc_videosoc_sdram_inti_p1_rddata_en = (soc_videosoc_sdram_phaseinjector1_command_issue_re & soc_videosoc_sdram_phaseinjector1_command_storage[5]);
assign soc_videosoc_sdram_inti_p1_wrdata = soc_videosoc_sdram_phaseinjector1_wrdata_storage;
assign soc_videosoc_sdram_inti_p1_wrdata_mask = 1'd0;
always @(*) begin
	soc_videosoc_sdram_inti_p2_cs_n <= 1'd1;
	soc_videosoc_sdram_inti_p2_ras_n <= 1'd1;
	soc_videosoc_sdram_inti_p2_we_n <= 1'd1;
	soc_videosoc_sdram_inti_p2_cas_n <= 1'd1;
	if (soc_videosoc_sdram_phaseinjector2_command_issue_re) begin
		soc_videosoc_sdram_inti_p2_cs_n <= (~soc_videosoc_sdram_phaseinjector2_command_storage[0]);
		soc_videosoc_sdram_inti_p2_we_n <= (~soc_videosoc_sdram_phaseinjector2_command_storage[1]);
		soc_videosoc_sdram_inti_p2_cas_n <= (~soc_videosoc_sdram_phaseinjector2_command_storage[2]);
		soc_videosoc_sdram_inti_p2_ras_n <= (~soc_videosoc_sdram_phaseinjector2_command_storage[3]);
	end else begin
		soc_videosoc_sdram_inti_p2_cs_n <= 1'd1;
		soc_videosoc_sdram_inti_p2_we_n <= 1'd1;
		soc_videosoc_sdram_inti_p2_cas_n <= 1'd1;
		soc_videosoc_sdram_inti_p2_ras_n <= 1'd1;
	end
end
assign soc_videosoc_sdram_inti_p2_address = soc_videosoc_sdram_phaseinjector2_address_storage;
assign soc_videosoc_sdram_inti_p2_bank = soc_videosoc_sdram_phaseinjector2_baddress_storage;
assign soc_videosoc_sdram_inti_p2_wrdata_en = (soc_videosoc_sdram_phaseinjector2_command_issue_re & soc_videosoc_sdram_phaseinjector2_command_storage[4]);
assign soc_videosoc_sdram_inti_p2_rddata_en = (soc_videosoc_sdram_phaseinjector2_command_issue_re & soc_videosoc_sdram_phaseinjector2_command_storage[5]);
assign soc_videosoc_sdram_inti_p2_wrdata = soc_videosoc_sdram_phaseinjector2_wrdata_storage;
assign soc_videosoc_sdram_inti_p2_wrdata_mask = 1'd0;
always @(*) begin
	soc_videosoc_sdram_inti_p3_ras_n <= 1'd1;
	soc_videosoc_sdram_inti_p3_we_n <= 1'd1;
	soc_videosoc_sdram_inti_p3_cas_n <= 1'd1;
	soc_videosoc_sdram_inti_p3_cs_n <= 1'd1;
	if (soc_videosoc_sdram_phaseinjector3_command_issue_re) begin
		soc_videosoc_sdram_inti_p3_cs_n <= (~soc_videosoc_sdram_phaseinjector3_command_storage[0]);
		soc_videosoc_sdram_inti_p3_we_n <= (~soc_videosoc_sdram_phaseinjector3_command_storage[1]);
		soc_videosoc_sdram_inti_p3_cas_n <= (~soc_videosoc_sdram_phaseinjector3_command_storage[2]);
		soc_videosoc_sdram_inti_p3_ras_n <= (~soc_videosoc_sdram_phaseinjector3_command_storage[3]);
	end else begin
		soc_videosoc_sdram_inti_p3_cs_n <= 1'd1;
		soc_videosoc_sdram_inti_p3_we_n <= 1'd1;
		soc_videosoc_sdram_inti_p3_cas_n <= 1'd1;
		soc_videosoc_sdram_inti_p3_ras_n <= 1'd1;
	end
end
assign soc_videosoc_sdram_inti_p3_address = soc_videosoc_sdram_phaseinjector3_address_storage;
assign soc_videosoc_sdram_inti_p3_bank = soc_videosoc_sdram_phaseinjector3_baddress_storage;
assign soc_videosoc_sdram_inti_p3_wrdata_en = (soc_videosoc_sdram_phaseinjector3_command_issue_re & soc_videosoc_sdram_phaseinjector3_command_storage[4]);
assign soc_videosoc_sdram_inti_p3_rddata_en = (soc_videosoc_sdram_phaseinjector3_command_issue_re & soc_videosoc_sdram_phaseinjector3_command_storage[5]);
assign soc_videosoc_sdram_inti_p3_wrdata = soc_videosoc_sdram_phaseinjector3_wrdata_storage;
assign soc_videosoc_sdram_inti_p3_wrdata_mask = 1'd0;
assign soc_videosoc_sdram_bankmachine0_req_valid = soc_videosoc_sdram_interface_bank0_valid;
assign soc_videosoc_sdram_interface_bank0_ready = soc_videosoc_sdram_bankmachine0_req_ready;
assign soc_videosoc_sdram_bankmachine0_req_we = soc_videosoc_sdram_interface_bank0_we;
assign soc_videosoc_sdram_bankmachine0_req_adr = soc_videosoc_sdram_interface_bank0_adr;
assign soc_videosoc_sdram_interface_bank0_lock = soc_videosoc_sdram_bankmachine0_req_lock;
assign soc_videosoc_sdram_interface_bank0_wdata_ready = soc_videosoc_sdram_bankmachine0_req_wdata_ready;
assign soc_videosoc_sdram_interface_bank0_rdata_valid = soc_videosoc_sdram_bankmachine0_req_rdata_valid;
assign soc_videosoc_sdram_bankmachine1_req_valid = soc_videosoc_sdram_interface_bank1_valid;
assign soc_videosoc_sdram_interface_bank1_ready = soc_videosoc_sdram_bankmachine1_req_ready;
assign soc_videosoc_sdram_bankmachine1_req_we = soc_videosoc_sdram_interface_bank1_we;
assign soc_videosoc_sdram_bankmachine1_req_adr = soc_videosoc_sdram_interface_bank1_adr;
assign soc_videosoc_sdram_interface_bank1_lock = soc_videosoc_sdram_bankmachine1_req_lock;
assign soc_videosoc_sdram_interface_bank1_wdata_ready = soc_videosoc_sdram_bankmachine1_req_wdata_ready;
assign soc_videosoc_sdram_interface_bank1_rdata_valid = soc_videosoc_sdram_bankmachine1_req_rdata_valid;
assign soc_videosoc_sdram_bankmachine2_req_valid = soc_videosoc_sdram_interface_bank2_valid;
assign soc_videosoc_sdram_interface_bank2_ready = soc_videosoc_sdram_bankmachine2_req_ready;
assign soc_videosoc_sdram_bankmachine2_req_we = soc_videosoc_sdram_interface_bank2_we;
assign soc_videosoc_sdram_bankmachine2_req_adr = soc_videosoc_sdram_interface_bank2_adr;
assign soc_videosoc_sdram_interface_bank2_lock = soc_videosoc_sdram_bankmachine2_req_lock;
assign soc_videosoc_sdram_interface_bank2_wdata_ready = soc_videosoc_sdram_bankmachine2_req_wdata_ready;
assign soc_videosoc_sdram_interface_bank2_rdata_valid = soc_videosoc_sdram_bankmachine2_req_rdata_valid;
assign soc_videosoc_sdram_bankmachine3_req_valid = soc_videosoc_sdram_interface_bank3_valid;
assign soc_videosoc_sdram_interface_bank3_ready = soc_videosoc_sdram_bankmachine3_req_ready;
assign soc_videosoc_sdram_bankmachine3_req_we = soc_videosoc_sdram_interface_bank3_we;
assign soc_videosoc_sdram_bankmachine3_req_adr = soc_videosoc_sdram_interface_bank3_adr;
assign soc_videosoc_sdram_interface_bank3_lock = soc_videosoc_sdram_bankmachine3_req_lock;
assign soc_videosoc_sdram_interface_bank3_wdata_ready = soc_videosoc_sdram_bankmachine3_req_wdata_ready;
assign soc_videosoc_sdram_interface_bank3_rdata_valid = soc_videosoc_sdram_bankmachine3_req_rdata_valid;
assign soc_videosoc_sdram_bankmachine4_req_valid = soc_videosoc_sdram_interface_bank4_valid;
assign soc_videosoc_sdram_interface_bank4_ready = soc_videosoc_sdram_bankmachine4_req_ready;
assign soc_videosoc_sdram_bankmachine4_req_we = soc_videosoc_sdram_interface_bank4_we;
assign soc_videosoc_sdram_bankmachine4_req_adr = soc_videosoc_sdram_interface_bank4_adr;
assign soc_videosoc_sdram_interface_bank4_lock = soc_videosoc_sdram_bankmachine4_req_lock;
assign soc_videosoc_sdram_interface_bank4_wdata_ready = soc_videosoc_sdram_bankmachine4_req_wdata_ready;
assign soc_videosoc_sdram_interface_bank4_rdata_valid = soc_videosoc_sdram_bankmachine4_req_rdata_valid;
assign soc_videosoc_sdram_bankmachine5_req_valid = soc_videosoc_sdram_interface_bank5_valid;
assign soc_videosoc_sdram_interface_bank5_ready = soc_videosoc_sdram_bankmachine5_req_ready;
assign soc_videosoc_sdram_bankmachine5_req_we = soc_videosoc_sdram_interface_bank5_we;
assign soc_videosoc_sdram_bankmachine5_req_adr = soc_videosoc_sdram_interface_bank5_adr;
assign soc_videosoc_sdram_interface_bank5_lock = soc_videosoc_sdram_bankmachine5_req_lock;
assign soc_videosoc_sdram_interface_bank5_wdata_ready = soc_videosoc_sdram_bankmachine5_req_wdata_ready;
assign soc_videosoc_sdram_interface_bank5_rdata_valid = soc_videosoc_sdram_bankmachine5_req_rdata_valid;
assign soc_videosoc_sdram_bankmachine6_req_valid = soc_videosoc_sdram_interface_bank6_valid;
assign soc_videosoc_sdram_interface_bank6_ready = soc_videosoc_sdram_bankmachine6_req_ready;
assign soc_videosoc_sdram_bankmachine6_req_we = soc_videosoc_sdram_interface_bank6_we;
assign soc_videosoc_sdram_bankmachine6_req_adr = soc_videosoc_sdram_interface_bank6_adr;
assign soc_videosoc_sdram_interface_bank6_lock = soc_videosoc_sdram_bankmachine6_req_lock;
assign soc_videosoc_sdram_interface_bank6_wdata_ready = soc_videosoc_sdram_bankmachine6_req_wdata_ready;
assign soc_videosoc_sdram_interface_bank6_rdata_valid = soc_videosoc_sdram_bankmachine6_req_rdata_valid;
assign soc_videosoc_sdram_bankmachine7_req_valid = soc_videosoc_sdram_interface_bank7_valid;
assign soc_videosoc_sdram_interface_bank7_ready = soc_videosoc_sdram_bankmachine7_req_ready;
assign soc_videosoc_sdram_bankmachine7_req_we = soc_videosoc_sdram_interface_bank7_we;
assign soc_videosoc_sdram_bankmachine7_req_adr = soc_videosoc_sdram_interface_bank7_adr;
assign soc_videosoc_sdram_interface_bank7_lock = soc_videosoc_sdram_bankmachine7_req_lock;
assign soc_videosoc_sdram_interface_bank7_wdata_ready = soc_videosoc_sdram_bankmachine7_req_wdata_ready;
assign soc_videosoc_sdram_interface_bank7_rdata_valid = soc_videosoc_sdram_bankmachine7_req_rdata_valid;
assign soc_videosoc_sdram_wait = (1'd1 & (~soc_videosoc_sdram_done));
assign soc_videosoc_sdram_done = (soc_videosoc_sdram_count == 1'd0);
always @(*) begin
	soc_videosoc_sdram_cmd_last <= 1'd0;
	soc_videosoc_sdram_seq_start <= 1'd0;
	soc_videosoc_sdram_cmd_valid <= 1'd0;
	vns_refresher_next_state <= 2'd0;
	vns_refresher_next_state <= vns_refresher_state;
	case (vns_refresher_state)
		1'd1: begin
			soc_videosoc_sdram_cmd_valid <= 1'd1;
			if (soc_videosoc_sdram_cmd_ready) begin
				soc_videosoc_sdram_seq_start <= 1'd1;
				vns_refresher_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if (soc_videosoc_sdram_seq_done) begin
				soc_videosoc_sdram_cmd_last <= 1'd1;
				vns_refresher_next_state <= 1'd0;
			end else begin
				soc_videosoc_sdram_cmd_valid <= 1'd1;
			end
		end
		default: begin
			if (soc_videosoc_sdram_done) begin
				vns_refresher_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videosoc_sdram_bankmachine0_sink_valid = soc_videosoc_sdram_bankmachine0_req_valid;
assign soc_videosoc_sdram_bankmachine0_req_ready = soc_videosoc_sdram_bankmachine0_sink_ready;
assign soc_videosoc_sdram_bankmachine0_sink_payload_we = soc_videosoc_sdram_bankmachine0_req_we;
assign soc_videosoc_sdram_bankmachine0_sink_payload_adr = soc_videosoc_sdram_bankmachine0_req_adr;
assign soc_videosoc_sdram_bankmachine0_source_ready = (soc_videosoc_sdram_bankmachine0_req_wdata_ready | soc_videosoc_sdram_bankmachine0_req_rdata_valid);
assign soc_videosoc_sdram_bankmachine0_req_lock = soc_videosoc_sdram_bankmachine0_source_valid;
assign soc_videosoc_sdram_bankmachine0_hit = (soc_videosoc_sdram_bankmachine0_openrow == soc_videosoc_sdram_bankmachine0_source_payload_adr[21:7]);
assign soc_videosoc_sdram_bankmachine0_cmd_payload_ba = 1'd0;
always @(*) begin
	soc_videosoc_sdram_bankmachine0_cmd_payload_a <= 15'd0;
	if (soc_videosoc_sdram_bankmachine0_sel_row_adr) begin
		soc_videosoc_sdram_bankmachine0_cmd_payload_a <= soc_videosoc_sdram_bankmachine0_source_payload_adr[21:7];
	end else begin
		soc_videosoc_sdram_bankmachine0_cmd_payload_a <= {soc_videosoc_sdram_bankmachine0_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign soc_videosoc_sdram_bankmachine0_wait = (~((soc_videosoc_sdram_bankmachine0_cmd_valid & soc_videosoc_sdram_bankmachine0_cmd_ready) & soc_videosoc_sdram_bankmachine0_cmd_payload_is_write));
assign soc_videosoc_sdram_bankmachine0_syncfifo0_din = {soc_videosoc_sdram_bankmachine0_fifo_in_last, soc_videosoc_sdram_bankmachine0_fifo_in_first, soc_videosoc_sdram_bankmachine0_fifo_in_payload_adr, soc_videosoc_sdram_bankmachine0_fifo_in_payload_we};
assign {soc_videosoc_sdram_bankmachine0_fifo_out_last, soc_videosoc_sdram_bankmachine0_fifo_out_first, soc_videosoc_sdram_bankmachine0_fifo_out_payload_adr, soc_videosoc_sdram_bankmachine0_fifo_out_payload_we} = soc_videosoc_sdram_bankmachine0_syncfifo0_dout;
assign soc_videosoc_sdram_bankmachine0_sink_ready = soc_videosoc_sdram_bankmachine0_syncfifo0_writable;
assign soc_videosoc_sdram_bankmachine0_syncfifo0_we = soc_videosoc_sdram_bankmachine0_sink_valid;
assign soc_videosoc_sdram_bankmachine0_fifo_in_first = soc_videosoc_sdram_bankmachine0_sink_first;
assign soc_videosoc_sdram_bankmachine0_fifo_in_last = soc_videosoc_sdram_bankmachine0_sink_last;
assign soc_videosoc_sdram_bankmachine0_fifo_in_payload_we = soc_videosoc_sdram_bankmachine0_sink_payload_we;
assign soc_videosoc_sdram_bankmachine0_fifo_in_payload_adr = soc_videosoc_sdram_bankmachine0_sink_payload_adr;
assign soc_videosoc_sdram_bankmachine0_source_valid = soc_videosoc_sdram_bankmachine0_syncfifo0_readable;
assign soc_videosoc_sdram_bankmachine0_source_first = soc_videosoc_sdram_bankmachine0_fifo_out_first;
assign soc_videosoc_sdram_bankmachine0_source_last = soc_videosoc_sdram_bankmachine0_fifo_out_last;
assign soc_videosoc_sdram_bankmachine0_source_payload_we = soc_videosoc_sdram_bankmachine0_fifo_out_payload_we;
assign soc_videosoc_sdram_bankmachine0_source_payload_adr = soc_videosoc_sdram_bankmachine0_fifo_out_payload_adr;
assign soc_videosoc_sdram_bankmachine0_syncfifo0_re = soc_videosoc_sdram_bankmachine0_source_ready;
always @(*) begin
	soc_videosoc_sdram_bankmachine0_wrport_adr <= 3'd0;
	if (soc_videosoc_sdram_bankmachine0_replace) begin
		soc_videosoc_sdram_bankmachine0_wrport_adr <= (soc_videosoc_sdram_bankmachine0_produce - 1'd1);
	end else begin
		soc_videosoc_sdram_bankmachine0_wrport_adr <= soc_videosoc_sdram_bankmachine0_produce;
	end
end
assign soc_videosoc_sdram_bankmachine0_wrport_dat_w = soc_videosoc_sdram_bankmachine0_syncfifo0_din;
assign soc_videosoc_sdram_bankmachine0_wrport_we = (soc_videosoc_sdram_bankmachine0_syncfifo0_we & (soc_videosoc_sdram_bankmachine0_syncfifo0_writable | soc_videosoc_sdram_bankmachine0_replace));
assign soc_videosoc_sdram_bankmachine0_do_read = (soc_videosoc_sdram_bankmachine0_syncfifo0_readable & soc_videosoc_sdram_bankmachine0_syncfifo0_re);
assign soc_videosoc_sdram_bankmachine0_rdport_adr = soc_videosoc_sdram_bankmachine0_consume;
assign soc_videosoc_sdram_bankmachine0_syncfifo0_dout = soc_videosoc_sdram_bankmachine0_rdport_dat_r;
assign soc_videosoc_sdram_bankmachine0_syncfifo0_writable = (soc_videosoc_sdram_bankmachine0_level != 4'd8);
assign soc_videosoc_sdram_bankmachine0_syncfifo0_readable = (soc_videosoc_sdram_bankmachine0_level != 1'd0);
assign soc_videosoc_sdram_bankmachine0_done = (soc_videosoc_sdram_bankmachine0_count == 1'd0);
always @(*) begin
	soc_videosoc_sdram_bankmachine0_track_open <= 1'd0;
	soc_videosoc_sdram_bankmachine0_track_close <= 1'd0;
	soc_videosoc_sdram_bankmachine0_cmd_payload_cas <= 1'd0;
	soc_videosoc_sdram_bankmachine0_cmd_payload_ras <= 1'd0;
	soc_videosoc_sdram_bankmachine0_cmd_payload_we <= 1'd0;
	soc_videosoc_sdram_bankmachine0_sel_row_adr <= 1'd0;
	soc_videosoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd0;
	soc_videosoc_sdram_bankmachine0_cmd_payload_is_read <= 1'd0;
	soc_videosoc_sdram_bankmachine0_cmd_payload_is_write <= 1'd0;
	soc_videosoc_sdram_bankmachine0_req_wdata_ready <= 1'd0;
	soc_videosoc_sdram_bankmachine0_req_rdata_valid <= 1'd0;
	vns_bankmachine0_next_state <= 3'd0;
	soc_videosoc_sdram_bankmachine0_refresh_gnt <= 1'd0;
	soc_videosoc_sdram_bankmachine0_cmd_valid <= 1'd0;
	vns_bankmachine0_next_state <= vns_bankmachine0_state;
	case (vns_bankmachine0_state)
		1'd1: begin
			if (soc_videosoc_sdram_bankmachine0_done) begin
				soc_videosoc_sdram_bankmachine0_cmd_valid <= 1'd1;
				if (soc_videosoc_sdram_bankmachine0_cmd_ready) begin
					vns_bankmachine0_next_state <= 3'd4;
				end
				soc_videosoc_sdram_bankmachine0_cmd_payload_ras <= 1'd1;
				soc_videosoc_sdram_bankmachine0_cmd_payload_we <= 1'd1;
				soc_videosoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine0_track_close <= 1'd1;
		end
		2'd2: begin
			soc_videosoc_sdram_bankmachine0_sel_row_adr <= 1'd1;
			soc_videosoc_sdram_bankmachine0_track_open <= 1'd1;
			soc_videosoc_sdram_bankmachine0_cmd_valid <= 1'd1;
			soc_videosoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd1;
			if (soc_videosoc_sdram_bankmachine0_cmd_ready) begin
				vns_bankmachine0_next_state <= 3'd6;
			end
			soc_videosoc_sdram_bankmachine0_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (soc_videosoc_sdram_bankmachine0_done) begin
				soc_videosoc_sdram_bankmachine0_refresh_gnt <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine0_track_close <= 1'd1;
			soc_videosoc_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videosoc_sdram_bankmachine0_refresh_req)) begin
				vns_bankmachine0_next_state <= 1'd0;
			end
		end
		3'd4: begin
			vns_bankmachine0_next_state <= 3'd5;
		end
		3'd5: begin
			vns_bankmachine0_next_state <= 2'd2;
		end
		3'd6: begin
			vns_bankmachine0_next_state <= 3'd7;
		end
		3'd7: begin
			vns_bankmachine0_next_state <= 1'd0;
		end
		default: begin
			if (soc_videosoc_sdram_bankmachine0_refresh_req) begin
				vns_bankmachine0_next_state <= 2'd3;
			end else begin
				if (soc_videosoc_sdram_bankmachine0_source_valid) begin
					if (soc_videosoc_sdram_bankmachine0_has_openrow) begin
						if (soc_videosoc_sdram_bankmachine0_hit) begin
							soc_videosoc_sdram_bankmachine0_cmd_valid <= 1'd1;
							if (soc_videosoc_sdram_bankmachine0_source_payload_we) begin
								soc_videosoc_sdram_bankmachine0_req_wdata_ready <= soc_videosoc_sdram_bankmachine0_cmd_ready;
								soc_videosoc_sdram_bankmachine0_cmd_payload_is_write <= 1'd1;
								soc_videosoc_sdram_bankmachine0_cmd_payload_we <= 1'd1;
							end else begin
								soc_videosoc_sdram_bankmachine0_req_rdata_valid <= soc_videosoc_sdram_bankmachine0_cmd_ready;
								soc_videosoc_sdram_bankmachine0_cmd_payload_is_read <= 1'd1;
							end
							soc_videosoc_sdram_bankmachine0_cmd_payload_cas <= 1'd1;
						end else begin
							vns_bankmachine0_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine0_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign soc_videosoc_sdram_bankmachine1_sink_valid = soc_videosoc_sdram_bankmachine1_req_valid;
assign soc_videosoc_sdram_bankmachine1_req_ready = soc_videosoc_sdram_bankmachine1_sink_ready;
assign soc_videosoc_sdram_bankmachine1_sink_payload_we = soc_videosoc_sdram_bankmachine1_req_we;
assign soc_videosoc_sdram_bankmachine1_sink_payload_adr = soc_videosoc_sdram_bankmachine1_req_adr;
assign soc_videosoc_sdram_bankmachine1_source_ready = (soc_videosoc_sdram_bankmachine1_req_wdata_ready | soc_videosoc_sdram_bankmachine1_req_rdata_valid);
assign soc_videosoc_sdram_bankmachine1_req_lock = soc_videosoc_sdram_bankmachine1_source_valid;
assign soc_videosoc_sdram_bankmachine1_hit = (soc_videosoc_sdram_bankmachine1_openrow == soc_videosoc_sdram_bankmachine1_source_payload_adr[21:7]);
assign soc_videosoc_sdram_bankmachine1_cmd_payload_ba = 1'd1;
always @(*) begin
	soc_videosoc_sdram_bankmachine1_cmd_payload_a <= 15'd0;
	if (soc_videosoc_sdram_bankmachine1_sel_row_adr) begin
		soc_videosoc_sdram_bankmachine1_cmd_payload_a <= soc_videosoc_sdram_bankmachine1_source_payload_adr[21:7];
	end else begin
		soc_videosoc_sdram_bankmachine1_cmd_payload_a <= {soc_videosoc_sdram_bankmachine1_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign soc_videosoc_sdram_bankmachine1_wait = (~((soc_videosoc_sdram_bankmachine1_cmd_valid & soc_videosoc_sdram_bankmachine1_cmd_ready) & soc_videosoc_sdram_bankmachine1_cmd_payload_is_write));
assign soc_videosoc_sdram_bankmachine1_syncfifo1_din = {soc_videosoc_sdram_bankmachine1_fifo_in_last, soc_videosoc_sdram_bankmachine1_fifo_in_first, soc_videosoc_sdram_bankmachine1_fifo_in_payload_adr, soc_videosoc_sdram_bankmachine1_fifo_in_payload_we};
assign {soc_videosoc_sdram_bankmachine1_fifo_out_last, soc_videosoc_sdram_bankmachine1_fifo_out_first, soc_videosoc_sdram_bankmachine1_fifo_out_payload_adr, soc_videosoc_sdram_bankmachine1_fifo_out_payload_we} = soc_videosoc_sdram_bankmachine1_syncfifo1_dout;
assign soc_videosoc_sdram_bankmachine1_sink_ready = soc_videosoc_sdram_bankmachine1_syncfifo1_writable;
assign soc_videosoc_sdram_bankmachine1_syncfifo1_we = soc_videosoc_sdram_bankmachine1_sink_valid;
assign soc_videosoc_sdram_bankmachine1_fifo_in_first = soc_videosoc_sdram_bankmachine1_sink_first;
assign soc_videosoc_sdram_bankmachine1_fifo_in_last = soc_videosoc_sdram_bankmachine1_sink_last;
assign soc_videosoc_sdram_bankmachine1_fifo_in_payload_we = soc_videosoc_sdram_bankmachine1_sink_payload_we;
assign soc_videosoc_sdram_bankmachine1_fifo_in_payload_adr = soc_videosoc_sdram_bankmachine1_sink_payload_adr;
assign soc_videosoc_sdram_bankmachine1_source_valid = soc_videosoc_sdram_bankmachine1_syncfifo1_readable;
assign soc_videosoc_sdram_bankmachine1_source_first = soc_videosoc_sdram_bankmachine1_fifo_out_first;
assign soc_videosoc_sdram_bankmachine1_source_last = soc_videosoc_sdram_bankmachine1_fifo_out_last;
assign soc_videosoc_sdram_bankmachine1_source_payload_we = soc_videosoc_sdram_bankmachine1_fifo_out_payload_we;
assign soc_videosoc_sdram_bankmachine1_source_payload_adr = soc_videosoc_sdram_bankmachine1_fifo_out_payload_adr;
assign soc_videosoc_sdram_bankmachine1_syncfifo1_re = soc_videosoc_sdram_bankmachine1_source_ready;
always @(*) begin
	soc_videosoc_sdram_bankmachine1_wrport_adr <= 3'd0;
	if (soc_videosoc_sdram_bankmachine1_replace) begin
		soc_videosoc_sdram_bankmachine1_wrport_adr <= (soc_videosoc_sdram_bankmachine1_produce - 1'd1);
	end else begin
		soc_videosoc_sdram_bankmachine1_wrport_adr <= soc_videosoc_sdram_bankmachine1_produce;
	end
end
assign soc_videosoc_sdram_bankmachine1_wrport_dat_w = soc_videosoc_sdram_bankmachine1_syncfifo1_din;
assign soc_videosoc_sdram_bankmachine1_wrport_we = (soc_videosoc_sdram_bankmachine1_syncfifo1_we & (soc_videosoc_sdram_bankmachine1_syncfifo1_writable | soc_videosoc_sdram_bankmachine1_replace));
assign soc_videosoc_sdram_bankmachine1_do_read = (soc_videosoc_sdram_bankmachine1_syncfifo1_readable & soc_videosoc_sdram_bankmachine1_syncfifo1_re);
assign soc_videosoc_sdram_bankmachine1_rdport_adr = soc_videosoc_sdram_bankmachine1_consume;
assign soc_videosoc_sdram_bankmachine1_syncfifo1_dout = soc_videosoc_sdram_bankmachine1_rdport_dat_r;
assign soc_videosoc_sdram_bankmachine1_syncfifo1_writable = (soc_videosoc_sdram_bankmachine1_level != 4'd8);
assign soc_videosoc_sdram_bankmachine1_syncfifo1_readable = (soc_videosoc_sdram_bankmachine1_level != 1'd0);
assign soc_videosoc_sdram_bankmachine1_done = (soc_videosoc_sdram_bankmachine1_count == 1'd0);
always @(*) begin
	soc_videosoc_sdram_bankmachine1_req_wdata_ready <= 1'd0;
	soc_videosoc_sdram_bankmachine1_req_rdata_valid <= 1'd0;
	soc_videosoc_sdram_bankmachine1_refresh_gnt <= 1'd0;
	soc_videosoc_sdram_bankmachine1_cmd_valid <= 1'd0;
	soc_videosoc_sdram_bankmachine1_track_open <= 1'd0;
	soc_videosoc_sdram_bankmachine1_track_close <= 1'd0;
	vns_bankmachine1_next_state <= 3'd0;
	soc_videosoc_sdram_bankmachine1_cmd_payload_ras <= 1'd0;
	soc_videosoc_sdram_bankmachine1_cmd_payload_cas <= 1'd0;
	soc_videosoc_sdram_bankmachine1_cmd_payload_we <= 1'd0;
	soc_videosoc_sdram_bankmachine1_sel_row_adr <= 1'd0;
	soc_videosoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd0;
	soc_videosoc_sdram_bankmachine1_cmd_payload_is_read <= 1'd0;
	soc_videosoc_sdram_bankmachine1_cmd_payload_is_write <= 1'd0;
	vns_bankmachine1_next_state <= vns_bankmachine1_state;
	case (vns_bankmachine1_state)
		1'd1: begin
			if (soc_videosoc_sdram_bankmachine1_done) begin
				soc_videosoc_sdram_bankmachine1_cmd_valid <= 1'd1;
				if (soc_videosoc_sdram_bankmachine1_cmd_ready) begin
					vns_bankmachine1_next_state <= 3'd4;
				end
				soc_videosoc_sdram_bankmachine1_cmd_payload_ras <= 1'd1;
				soc_videosoc_sdram_bankmachine1_cmd_payload_we <= 1'd1;
				soc_videosoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine1_track_close <= 1'd1;
		end
		2'd2: begin
			soc_videosoc_sdram_bankmachine1_sel_row_adr <= 1'd1;
			soc_videosoc_sdram_bankmachine1_track_open <= 1'd1;
			soc_videosoc_sdram_bankmachine1_cmd_valid <= 1'd1;
			soc_videosoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd1;
			if (soc_videosoc_sdram_bankmachine1_cmd_ready) begin
				vns_bankmachine1_next_state <= 3'd6;
			end
			soc_videosoc_sdram_bankmachine1_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (soc_videosoc_sdram_bankmachine1_done) begin
				soc_videosoc_sdram_bankmachine1_refresh_gnt <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine1_track_close <= 1'd1;
			soc_videosoc_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videosoc_sdram_bankmachine1_refresh_req)) begin
				vns_bankmachine1_next_state <= 1'd0;
			end
		end
		3'd4: begin
			vns_bankmachine1_next_state <= 3'd5;
		end
		3'd5: begin
			vns_bankmachine1_next_state <= 2'd2;
		end
		3'd6: begin
			vns_bankmachine1_next_state <= 3'd7;
		end
		3'd7: begin
			vns_bankmachine1_next_state <= 1'd0;
		end
		default: begin
			if (soc_videosoc_sdram_bankmachine1_refresh_req) begin
				vns_bankmachine1_next_state <= 2'd3;
			end else begin
				if (soc_videosoc_sdram_bankmachine1_source_valid) begin
					if (soc_videosoc_sdram_bankmachine1_has_openrow) begin
						if (soc_videosoc_sdram_bankmachine1_hit) begin
							soc_videosoc_sdram_bankmachine1_cmd_valid <= 1'd1;
							if (soc_videosoc_sdram_bankmachine1_source_payload_we) begin
								soc_videosoc_sdram_bankmachine1_req_wdata_ready <= soc_videosoc_sdram_bankmachine1_cmd_ready;
								soc_videosoc_sdram_bankmachine1_cmd_payload_is_write <= 1'd1;
								soc_videosoc_sdram_bankmachine1_cmd_payload_we <= 1'd1;
							end else begin
								soc_videosoc_sdram_bankmachine1_req_rdata_valid <= soc_videosoc_sdram_bankmachine1_cmd_ready;
								soc_videosoc_sdram_bankmachine1_cmd_payload_is_read <= 1'd1;
							end
							soc_videosoc_sdram_bankmachine1_cmd_payload_cas <= 1'd1;
						end else begin
							vns_bankmachine1_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine1_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign soc_videosoc_sdram_bankmachine2_sink_valid = soc_videosoc_sdram_bankmachine2_req_valid;
assign soc_videosoc_sdram_bankmachine2_req_ready = soc_videosoc_sdram_bankmachine2_sink_ready;
assign soc_videosoc_sdram_bankmachine2_sink_payload_we = soc_videosoc_sdram_bankmachine2_req_we;
assign soc_videosoc_sdram_bankmachine2_sink_payload_adr = soc_videosoc_sdram_bankmachine2_req_adr;
assign soc_videosoc_sdram_bankmachine2_source_ready = (soc_videosoc_sdram_bankmachine2_req_wdata_ready | soc_videosoc_sdram_bankmachine2_req_rdata_valid);
assign soc_videosoc_sdram_bankmachine2_req_lock = soc_videosoc_sdram_bankmachine2_source_valid;
assign soc_videosoc_sdram_bankmachine2_hit = (soc_videosoc_sdram_bankmachine2_openrow == soc_videosoc_sdram_bankmachine2_source_payload_adr[21:7]);
assign soc_videosoc_sdram_bankmachine2_cmd_payload_ba = 2'd2;
always @(*) begin
	soc_videosoc_sdram_bankmachine2_cmd_payload_a <= 15'd0;
	if (soc_videosoc_sdram_bankmachine2_sel_row_adr) begin
		soc_videosoc_sdram_bankmachine2_cmd_payload_a <= soc_videosoc_sdram_bankmachine2_source_payload_adr[21:7];
	end else begin
		soc_videosoc_sdram_bankmachine2_cmd_payload_a <= {soc_videosoc_sdram_bankmachine2_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign soc_videosoc_sdram_bankmachine2_wait = (~((soc_videosoc_sdram_bankmachine2_cmd_valid & soc_videosoc_sdram_bankmachine2_cmd_ready) & soc_videosoc_sdram_bankmachine2_cmd_payload_is_write));
assign soc_videosoc_sdram_bankmachine2_syncfifo2_din = {soc_videosoc_sdram_bankmachine2_fifo_in_last, soc_videosoc_sdram_bankmachine2_fifo_in_first, soc_videosoc_sdram_bankmachine2_fifo_in_payload_adr, soc_videosoc_sdram_bankmachine2_fifo_in_payload_we};
assign {soc_videosoc_sdram_bankmachine2_fifo_out_last, soc_videosoc_sdram_bankmachine2_fifo_out_first, soc_videosoc_sdram_bankmachine2_fifo_out_payload_adr, soc_videosoc_sdram_bankmachine2_fifo_out_payload_we} = soc_videosoc_sdram_bankmachine2_syncfifo2_dout;
assign soc_videosoc_sdram_bankmachine2_sink_ready = soc_videosoc_sdram_bankmachine2_syncfifo2_writable;
assign soc_videosoc_sdram_bankmachine2_syncfifo2_we = soc_videosoc_sdram_bankmachine2_sink_valid;
assign soc_videosoc_sdram_bankmachine2_fifo_in_first = soc_videosoc_sdram_bankmachine2_sink_first;
assign soc_videosoc_sdram_bankmachine2_fifo_in_last = soc_videosoc_sdram_bankmachine2_sink_last;
assign soc_videosoc_sdram_bankmachine2_fifo_in_payload_we = soc_videosoc_sdram_bankmachine2_sink_payload_we;
assign soc_videosoc_sdram_bankmachine2_fifo_in_payload_adr = soc_videosoc_sdram_bankmachine2_sink_payload_adr;
assign soc_videosoc_sdram_bankmachine2_source_valid = soc_videosoc_sdram_bankmachine2_syncfifo2_readable;
assign soc_videosoc_sdram_bankmachine2_source_first = soc_videosoc_sdram_bankmachine2_fifo_out_first;
assign soc_videosoc_sdram_bankmachine2_source_last = soc_videosoc_sdram_bankmachine2_fifo_out_last;
assign soc_videosoc_sdram_bankmachine2_source_payload_we = soc_videosoc_sdram_bankmachine2_fifo_out_payload_we;
assign soc_videosoc_sdram_bankmachine2_source_payload_adr = soc_videosoc_sdram_bankmachine2_fifo_out_payload_adr;
assign soc_videosoc_sdram_bankmachine2_syncfifo2_re = soc_videosoc_sdram_bankmachine2_source_ready;
always @(*) begin
	soc_videosoc_sdram_bankmachine2_wrport_adr <= 3'd0;
	if (soc_videosoc_sdram_bankmachine2_replace) begin
		soc_videosoc_sdram_bankmachine2_wrport_adr <= (soc_videosoc_sdram_bankmachine2_produce - 1'd1);
	end else begin
		soc_videosoc_sdram_bankmachine2_wrport_adr <= soc_videosoc_sdram_bankmachine2_produce;
	end
end
assign soc_videosoc_sdram_bankmachine2_wrport_dat_w = soc_videosoc_sdram_bankmachine2_syncfifo2_din;
assign soc_videosoc_sdram_bankmachine2_wrport_we = (soc_videosoc_sdram_bankmachine2_syncfifo2_we & (soc_videosoc_sdram_bankmachine2_syncfifo2_writable | soc_videosoc_sdram_bankmachine2_replace));
assign soc_videosoc_sdram_bankmachine2_do_read = (soc_videosoc_sdram_bankmachine2_syncfifo2_readable & soc_videosoc_sdram_bankmachine2_syncfifo2_re);
assign soc_videosoc_sdram_bankmachine2_rdport_adr = soc_videosoc_sdram_bankmachine2_consume;
assign soc_videosoc_sdram_bankmachine2_syncfifo2_dout = soc_videosoc_sdram_bankmachine2_rdport_dat_r;
assign soc_videosoc_sdram_bankmachine2_syncfifo2_writable = (soc_videosoc_sdram_bankmachine2_level != 4'd8);
assign soc_videosoc_sdram_bankmachine2_syncfifo2_readable = (soc_videosoc_sdram_bankmachine2_level != 1'd0);
assign soc_videosoc_sdram_bankmachine2_done = (soc_videosoc_sdram_bankmachine2_count == 1'd0);
always @(*) begin
	soc_videosoc_sdram_bankmachine2_track_close <= 1'd0;
	soc_videosoc_sdram_bankmachine2_cmd_payload_cas <= 1'd0;
	soc_videosoc_sdram_bankmachine2_cmd_payload_ras <= 1'd0;
	soc_videosoc_sdram_bankmachine2_cmd_payload_we <= 1'd0;
	soc_videosoc_sdram_bankmachine2_sel_row_adr <= 1'd0;
	soc_videosoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd0;
	soc_videosoc_sdram_bankmachine2_cmd_payload_is_read <= 1'd0;
	soc_videosoc_sdram_bankmachine2_cmd_payload_is_write <= 1'd0;
	soc_videosoc_sdram_bankmachine2_req_wdata_ready <= 1'd0;
	vns_bankmachine2_next_state <= 3'd0;
	soc_videosoc_sdram_bankmachine2_req_rdata_valid <= 1'd0;
	soc_videosoc_sdram_bankmachine2_refresh_gnt <= 1'd0;
	soc_videosoc_sdram_bankmachine2_cmd_valid <= 1'd0;
	soc_videosoc_sdram_bankmachine2_track_open <= 1'd0;
	vns_bankmachine2_next_state <= vns_bankmachine2_state;
	case (vns_bankmachine2_state)
		1'd1: begin
			if (soc_videosoc_sdram_bankmachine2_done) begin
				soc_videosoc_sdram_bankmachine2_cmd_valid <= 1'd1;
				if (soc_videosoc_sdram_bankmachine2_cmd_ready) begin
					vns_bankmachine2_next_state <= 3'd4;
				end
				soc_videosoc_sdram_bankmachine2_cmd_payload_ras <= 1'd1;
				soc_videosoc_sdram_bankmachine2_cmd_payload_we <= 1'd1;
				soc_videosoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine2_track_close <= 1'd1;
		end
		2'd2: begin
			soc_videosoc_sdram_bankmachine2_sel_row_adr <= 1'd1;
			soc_videosoc_sdram_bankmachine2_track_open <= 1'd1;
			soc_videosoc_sdram_bankmachine2_cmd_valid <= 1'd1;
			soc_videosoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd1;
			if (soc_videosoc_sdram_bankmachine2_cmd_ready) begin
				vns_bankmachine2_next_state <= 3'd6;
			end
			soc_videosoc_sdram_bankmachine2_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (soc_videosoc_sdram_bankmachine2_done) begin
				soc_videosoc_sdram_bankmachine2_refresh_gnt <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine2_track_close <= 1'd1;
			soc_videosoc_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videosoc_sdram_bankmachine2_refresh_req)) begin
				vns_bankmachine2_next_state <= 1'd0;
			end
		end
		3'd4: begin
			vns_bankmachine2_next_state <= 3'd5;
		end
		3'd5: begin
			vns_bankmachine2_next_state <= 2'd2;
		end
		3'd6: begin
			vns_bankmachine2_next_state <= 3'd7;
		end
		3'd7: begin
			vns_bankmachine2_next_state <= 1'd0;
		end
		default: begin
			if (soc_videosoc_sdram_bankmachine2_refresh_req) begin
				vns_bankmachine2_next_state <= 2'd3;
			end else begin
				if (soc_videosoc_sdram_bankmachine2_source_valid) begin
					if (soc_videosoc_sdram_bankmachine2_has_openrow) begin
						if (soc_videosoc_sdram_bankmachine2_hit) begin
							soc_videosoc_sdram_bankmachine2_cmd_valid <= 1'd1;
							if (soc_videosoc_sdram_bankmachine2_source_payload_we) begin
								soc_videosoc_sdram_bankmachine2_req_wdata_ready <= soc_videosoc_sdram_bankmachine2_cmd_ready;
								soc_videosoc_sdram_bankmachine2_cmd_payload_is_write <= 1'd1;
								soc_videosoc_sdram_bankmachine2_cmd_payload_we <= 1'd1;
							end else begin
								soc_videosoc_sdram_bankmachine2_req_rdata_valid <= soc_videosoc_sdram_bankmachine2_cmd_ready;
								soc_videosoc_sdram_bankmachine2_cmd_payload_is_read <= 1'd1;
							end
							soc_videosoc_sdram_bankmachine2_cmd_payload_cas <= 1'd1;
						end else begin
							vns_bankmachine2_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine2_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign soc_videosoc_sdram_bankmachine3_sink_valid = soc_videosoc_sdram_bankmachine3_req_valid;
assign soc_videosoc_sdram_bankmachine3_req_ready = soc_videosoc_sdram_bankmachine3_sink_ready;
assign soc_videosoc_sdram_bankmachine3_sink_payload_we = soc_videosoc_sdram_bankmachine3_req_we;
assign soc_videosoc_sdram_bankmachine3_sink_payload_adr = soc_videosoc_sdram_bankmachine3_req_adr;
assign soc_videosoc_sdram_bankmachine3_source_ready = (soc_videosoc_sdram_bankmachine3_req_wdata_ready | soc_videosoc_sdram_bankmachine3_req_rdata_valid);
assign soc_videosoc_sdram_bankmachine3_req_lock = soc_videosoc_sdram_bankmachine3_source_valid;
assign soc_videosoc_sdram_bankmachine3_hit = (soc_videosoc_sdram_bankmachine3_openrow == soc_videosoc_sdram_bankmachine3_source_payload_adr[21:7]);
assign soc_videosoc_sdram_bankmachine3_cmd_payload_ba = 2'd3;
always @(*) begin
	soc_videosoc_sdram_bankmachine3_cmd_payload_a <= 15'd0;
	if (soc_videosoc_sdram_bankmachine3_sel_row_adr) begin
		soc_videosoc_sdram_bankmachine3_cmd_payload_a <= soc_videosoc_sdram_bankmachine3_source_payload_adr[21:7];
	end else begin
		soc_videosoc_sdram_bankmachine3_cmd_payload_a <= {soc_videosoc_sdram_bankmachine3_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign soc_videosoc_sdram_bankmachine3_wait = (~((soc_videosoc_sdram_bankmachine3_cmd_valid & soc_videosoc_sdram_bankmachine3_cmd_ready) & soc_videosoc_sdram_bankmachine3_cmd_payload_is_write));
assign soc_videosoc_sdram_bankmachine3_syncfifo3_din = {soc_videosoc_sdram_bankmachine3_fifo_in_last, soc_videosoc_sdram_bankmachine3_fifo_in_first, soc_videosoc_sdram_bankmachine3_fifo_in_payload_adr, soc_videosoc_sdram_bankmachine3_fifo_in_payload_we};
assign {soc_videosoc_sdram_bankmachine3_fifo_out_last, soc_videosoc_sdram_bankmachine3_fifo_out_first, soc_videosoc_sdram_bankmachine3_fifo_out_payload_adr, soc_videosoc_sdram_bankmachine3_fifo_out_payload_we} = soc_videosoc_sdram_bankmachine3_syncfifo3_dout;
assign soc_videosoc_sdram_bankmachine3_sink_ready = soc_videosoc_sdram_bankmachine3_syncfifo3_writable;
assign soc_videosoc_sdram_bankmachine3_syncfifo3_we = soc_videosoc_sdram_bankmachine3_sink_valid;
assign soc_videosoc_sdram_bankmachine3_fifo_in_first = soc_videosoc_sdram_bankmachine3_sink_first;
assign soc_videosoc_sdram_bankmachine3_fifo_in_last = soc_videosoc_sdram_bankmachine3_sink_last;
assign soc_videosoc_sdram_bankmachine3_fifo_in_payload_we = soc_videosoc_sdram_bankmachine3_sink_payload_we;
assign soc_videosoc_sdram_bankmachine3_fifo_in_payload_adr = soc_videosoc_sdram_bankmachine3_sink_payload_adr;
assign soc_videosoc_sdram_bankmachine3_source_valid = soc_videosoc_sdram_bankmachine3_syncfifo3_readable;
assign soc_videosoc_sdram_bankmachine3_source_first = soc_videosoc_sdram_bankmachine3_fifo_out_first;
assign soc_videosoc_sdram_bankmachine3_source_last = soc_videosoc_sdram_bankmachine3_fifo_out_last;
assign soc_videosoc_sdram_bankmachine3_source_payload_we = soc_videosoc_sdram_bankmachine3_fifo_out_payload_we;
assign soc_videosoc_sdram_bankmachine3_source_payload_adr = soc_videosoc_sdram_bankmachine3_fifo_out_payload_adr;
assign soc_videosoc_sdram_bankmachine3_syncfifo3_re = soc_videosoc_sdram_bankmachine3_source_ready;
always @(*) begin
	soc_videosoc_sdram_bankmachine3_wrport_adr <= 3'd0;
	if (soc_videosoc_sdram_bankmachine3_replace) begin
		soc_videosoc_sdram_bankmachine3_wrport_adr <= (soc_videosoc_sdram_bankmachine3_produce - 1'd1);
	end else begin
		soc_videosoc_sdram_bankmachine3_wrport_adr <= soc_videosoc_sdram_bankmachine3_produce;
	end
end
assign soc_videosoc_sdram_bankmachine3_wrport_dat_w = soc_videosoc_sdram_bankmachine3_syncfifo3_din;
assign soc_videosoc_sdram_bankmachine3_wrport_we = (soc_videosoc_sdram_bankmachine3_syncfifo3_we & (soc_videosoc_sdram_bankmachine3_syncfifo3_writable | soc_videosoc_sdram_bankmachine3_replace));
assign soc_videosoc_sdram_bankmachine3_do_read = (soc_videosoc_sdram_bankmachine3_syncfifo3_readable & soc_videosoc_sdram_bankmachine3_syncfifo3_re);
assign soc_videosoc_sdram_bankmachine3_rdport_adr = soc_videosoc_sdram_bankmachine3_consume;
assign soc_videosoc_sdram_bankmachine3_syncfifo3_dout = soc_videosoc_sdram_bankmachine3_rdport_dat_r;
assign soc_videosoc_sdram_bankmachine3_syncfifo3_writable = (soc_videosoc_sdram_bankmachine3_level != 4'd8);
assign soc_videosoc_sdram_bankmachine3_syncfifo3_readable = (soc_videosoc_sdram_bankmachine3_level != 1'd0);
assign soc_videosoc_sdram_bankmachine3_done = (soc_videosoc_sdram_bankmachine3_count == 1'd0);
always @(*) begin
	soc_videosoc_sdram_bankmachine3_cmd_valid <= 1'd0;
	vns_bankmachine3_next_state <= 3'd0;
	soc_videosoc_sdram_bankmachine3_track_open <= 1'd0;
	soc_videosoc_sdram_bankmachine3_track_close <= 1'd0;
	soc_videosoc_sdram_bankmachine3_cmd_payload_cas <= 1'd0;
	soc_videosoc_sdram_bankmachine3_cmd_payload_ras <= 1'd0;
	soc_videosoc_sdram_bankmachine3_cmd_payload_we <= 1'd0;
	soc_videosoc_sdram_bankmachine3_sel_row_adr <= 1'd0;
	soc_videosoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd0;
	soc_videosoc_sdram_bankmachine3_cmd_payload_is_read <= 1'd0;
	soc_videosoc_sdram_bankmachine3_cmd_payload_is_write <= 1'd0;
	soc_videosoc_sdram_bankmachine3_req_wdata_ready <= 1'd0;
	soc_videosoc_sdram_bankmachine3_req_rdata_valid <= 1'd0;
	soc_videosoc_sdram_bankmachine3_refresh_gnt <= 1'd0;
	vns_bankmachine3_next_state <= vns_bankmachine3_state;
	case (vns_bankmachine3_state)
		1'd1: begin
			if (soc_videosoc_sdram_bankmachine3_done) begin
				soc_videosoc_sdram_bankmachine3_cmd_valid <= 1'd1;
				if (soc_videosoc_sdram_bankmachine3_cmd_ready) begin
					vns_bankmachine3_next_state <= 3'd4;
				end
				soc_videosoc_sdram_bankmachine3_cmd_payload_ras <= 1'd1;
				soc_videosoc_sdram_bankmachine3_cmd_payload_we <= 1'd1;
				soc_videosoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine3_track_close <= 1'd1;
		end
		2'd2: begin
			soc_videosoc_sdram_bankmachine3_sel_row_adr <= 1'd1;
			soc_videosoc_sdram_bankmachine3_track_open <= 1'd1;
			soc_videosoc_sdram_bankmachine3_cmd_valid <= 1'd1;
			soc_videosoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd1;
			if (soc_videosoc_sdram_bankmachine3_cmd_ready) begin
				vns_bankmachine3_next_state <= 3'd6;
			end
			soc_videosoc_sdram_bankmachine3_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (soc_videosoc_sdram_bankmachine3_done) begin
				soc_videosoc_sdram_bankmachine3_refresh_gnt <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine3_track_close <= 1'd1;
			soc_videosoc_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videosoc_sdram_bankmachine3_refresh_req)) begin
				vns_bankmachine3_next_state <= 1'd0;
			end
		end
		3'd4: begin
			vns_bankmachine3_next_state <= 3'd5;
		end
		3'd5: begin
			vns_bankmachine3_next_state <= 2'd2;
		end
		3'd6: begin
			vns_bankmachine3_next_state <= 3'd7;
		end
		3'd7: begin
			vns_bankmachine3_next_state <= 1'd0;
		end
		default: begin
			if (soc_videosoc_sdram_bankmachine3_refresh_req) begin
				vns_bankmachine3_next_state <= 2'd3;
			end else begin
				if (soc_videosoc_sdram_bankmachine3_source_valid) begin
					if (soc_videosoc_sdram_bankmachine3_has_openrow) begin
						if (soc_videosoc_sdram_bankmachine3_hit) begin
							soc_videosoc_sdram_bankmachine3_cmd_valid <= 1'd1;
							if (soc_videosoc_sdram_bankmachine3_source_payload_we) begin
								soc_videosoc_sdram_bankmachine3_req_wdata_ready <= soc_videosoc_sdram_bankmachine3_cmd_ready;
								soc_videosoc_sdram_bankmachine3_cmd_payload_is_write <= 1'd1;
								soc_videosoc_sdram_bankmachine3_cmd_payload_we <= 1'd1;
							end else begin
								soc_videosoc_sdram_bankmachine3_req_rdata_valid <= soc_videosoc_sdram_bankmachine3_cmd_ready;
								soc_videosoc_sdram_bankmachine3_cmd_payload_is_read <= 1'd1;
							end
							soc_videosoc_sdram_bankmachine3_cmd_payload_cas <= 1'd1;
						end else begin
							vns_bankmachine3_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine3_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign soc_videosoc_sdram_bankmachine4_sink_valid = soc_videosoc_sdram_bankmachine4_req_valid;
assign soc_videosoc_sdram_bankmachine4_req_ready = soc_videosoc_sdram_bankmachine4_sink_ready;
assign soc_videosoc_sdram_bankmachine4_sink_payload_we = soc_videosoc_sdram_bankmachine4_req_we;
assign soc_videosoc_sdram_bankmachine4_sink_payload_adr = soc_videosoc_sdram_bankmachine4_req_adr;
assign soc_videosoc_sdram_bankmachine4_source_ready = (soc_videosoc_sdram_bankmachine4_req_wdata_ready | soc_videosoc_sdram_bankmachine4_req_rdata_valid);
assign soc_videosoc_sdram_bankmachine4_req_lock = soc_videosoc_sdram_bankmachine4_source_valid;
assign soc_videosoc_sdram_bankmachine4_hit = (soc_videosoc_sdram_bankmachine4_openrow == soc_videosoc_sdram_bankmachine4_source_payload_adr[21:7]);
assign soc_videosoc_sdram_bankmachine4_cmd_payload_ba = 3'd4;
always @(*) begin
	soc_videosoc_sdram_bankmachine4_cmd_payload_a <= 15'd0;
	if (soc_videosoc_sdram_bankmachine4_sel_row_adr) begin
		soc_videosoc_sdram_bankmachine4_cmd_payload_a <= soc_videosoc_sdram_bankmachine4_source_payload_adr[21:7];
	end else begin
		soc_videosoc_sdram_bankmachine4_cmd_payload_a <= {soc_videosoc_sdram_bankmachine4_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign soc_videosoc_sdram_bankmachine4_wait = (~((soc_videosoc_sdram_bankmachine4_cmd_valid & soc_videosoc_sdram_bankmachine4_cmd_ready) & soc_videosoc_sdram_bankmachine4_cmd_payload_is_write));
assign soc_videosoc_sdram_bankmachine4_syncfifo4_din = {soc_videosoc_sdram_bankmachine4_fifo_in_last, soc_videosoc_sdram_bankmachine4_fifo_in_first, soc_videosoc_sdram_bankmachine4_fifo_in_payload_adr, soc_videosoc_sdram_bankmachine4_fifo_in_payload_we};
assign {soc_videosoc_sdram_bankmachine4_fifo_out_last, soc_videosoc_sdram_bankmachine4_fifo_out_first, soc_videosoc_sdram_bankmachine4_fifo_out_payload_adr, soc_videosoc_sdram_bankmachine4_fifo_out_payload_we} = soc_videosoc_sdram_bankmachine4_syncfifo4_dout;
assign soc_videosoc_sdram_bankmachine4_sink_ready = soc_videosoc_sdram_bankmachine4_syncfifo4_writable;
assign soc_videosoc_sdram_bankmachine4_syncfifo4_we = soc_videosoc_sdram_bankmachine4_sink_valid;
assign soc_videosoc_sdram_bankmachine4_fifo_in_first = soc_videosoc_sdram_bankmachine4_sink_first;
assign soc_videosoc_sdram_bankmachine4_fifo_in_last = soc_videosoc_sdram_bankmachine4_sink_last;
assign soc_videosoc_sdram_bankmachine4_fifo_in_payload_we = soc_videosoc_sdram_bankmachine4_sink_payload_we;
assign soc_videosoc_sdram_bankmachine4_fifo_in_payload_adr = soc_videosoc_sdram_bankmachine4_sink_payload_adr;
assign soc_videosoc_sdram_bankmachine4_source_valid = soc_videosoc_sdram_bankmachine4_syncfifo4_readable;
assign soc_videosoc_sdram_bankmachine4_source_first = soc_videosoc_sdram_bankmachine4_fifo_out_first;
assign soc_videosoc_sdram_bankmachine4_source_last = soc_videosoc_sdram_bankmachine4_fifo_out_last;
assign soc_videosoc_sdram_bankmachine4_source_payload_we = soc_videosoc_sdram_bankmachine4_fifo_out_payload_we;
assign soc_videosoc_sdram_bankmachine4_source_payload_adr = soc_videosoc_sdram_bankmachine4_fifo_out_payload_adr;
assign soc_videosoc_sdram_bankmachine4_syncfifo4_re = soc_videosoc_sdram_bankmachine4_source_ready;
always @(*) begin
	soc_videosoc_sdram_bankmachine4_wrport_adr <= 3'd0;
	if (soc_videosoc_sdram_bankmachine4_replace) begin
		soc_videosoc_sdram_bankmachine4_wrport_adr <= (soc_videosoc_sdram_bankmachine4_produce - 1'd1);
	end else begin
		soc_videosoc_sdram_bankmachine4_wrport_adr <= soc_videosoc_sdram_bankmachine4_produce;
	end
end
assign soc_videosoc_sdram_bankmachine4_wrport_dat_w = soc_videosoc_sdram_bankmachine4_syncfifo4_din;
assign soc_videosoc_sdram_bankmachine4_wrport_we = (soc_videosoc_sdram_bankmachine4_syncfifo4_we & (soc_videosoc_sdram_bankmachine4_syncfifo4_writable | soc_videosoc_sdram_bankmachine4_replace));
assign soc_videosoc_sdram_bankmachine4_do_read = (soc_videosoc_sdram_bankmachine4_syncfifo4_readable & soc_videosoc_sdram_bankmachine4_syncfifo4_re);
assign soc_videosoc_sdram_bankmachine4_rdport_adr = soc_videosoc_sdram_bankmachine4_consume;
assign soc_videosoc_sdram_bankmachine4_syncfifo4_dout = soc_videosoc_sdram_bankmachine4_rdport_dat_r;
assign soc_videosoc_sdram_bankmachine4_syncfifo4_writable = (soc_videosoc_sdram_bankmachine4_level != 4'd8);
assign soc_videosoc_sdram_bankmachine4_syncfifo4_readable = (soc_videosoc_sdram_bankmachine4_level != 1'd0);
assign soc_videosoc_sdram_bankmachine4_done = (soc_videosoc_sdram_bankmachine4_count == 1'd0);
always @(*) begin
	soc_videosoc_sdram_bankmachine4_cmd_payload_is_read <= 1'd0;
	vns_bankmachine4_next_state <= 3'd0;
	soc_videosoc_sdram_bankmachine4_cmd_payload_is_write <= 1'd0;
	soc_videosoc_sdram_bankmachine4_req_wdata_ready <= 1'd0;
	soc_videosoc_sdram_bankmachine4_req_rdata_valid <= 1'd0;
	soc_videosoc_sdram_bankmachine4_refresh_gnt <= 1'd0;
	soc_videosoc_sdram_bankmachine4_cmd_payload_cas <= 1'd0;
	soc_videosoc_sdram_bankmachine4_cmd_valid <= 1'd0;
	soc_videosoc_sdram_bankmachine4_track_open <= 1'd0;
	soc_videosoc_sdram_bankmachine4_track_close <= 1'd0;
	soc_videosoc_sdram_bankmachine4_cmd_payload_ras <= 1'd0;
	soc_videosoc_sdram_bankmachine4_cmd_payload_we <= 1'd0;
	soc_videosoc_sdram_bankmachine4_sel_row_adr <= 1'd0;
	soc_videosoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd0;
	vns_bankmachine4_next_state <= vns_bankmachine4_state;
	case (vns_bankmachine4_state)
		1'd1: begin
			if (soc_videosoc_sdram_bankmachine4_done) begin
				soc_videosoc_sdram_bankmachine4_cmd_valid <= 1'd1;
				if (soc_videosoc_sdram_bankmachine4_cmd_ready) begin
					vns_bankmachine4_next_state <= 3'd4;
				end
				soc_videosoc_sdram_bankmachine4_cmd_payload_ras <= 1'd1;
				soc_videosoc_sdram_bankmachine4_cmd_payload_we <= 1'd1;
				soc_videosoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine4_track_close <= 1'd1;
		end
		2'd2: begin
			soc_videosoc_sdram_bankmachine4_sel_row_adr <= 1'd1;
			soc_videosoc_sdram_bankmachine4_track_open <= 1'd1;
			soc_videosoc_sdram_bankmachine4_cmd_valid <= 1'd1;
			soc_videosoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd1;
			if (soc_videosoc_sdram_bankmachine4_cmd_ready) begin
				vns_bankmachine4_next_state <= 3'd6;
			end
			soc_videosoc_sdram_bankmachine4_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (soc_videosoc_sdram_bankmachine4_done) begin
				soc_videosoc_sdram_bankmachine4_refresh_gnt <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine4_track_close <= 1'd1;
			soc_videosoc_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videosoc_sdram_bankmachine4_refresh_req)) begin
				vns_bankmachine4_next_state <= 1'd0;
			end
		end
		3'd4: begin
			vns_bankmachine4_next_state <= 3'd5;
		end
		3'd5: begin
			vns_bankmachine4_next_state <= 2'd2;
		end
		3'd6: begin
			vns_bankmachine4_next_state <= 3'd7;
		end
		3'd7: begin
			vns_bankmachine4_next_state <= 1'd0;
		end
		default: begin
			if (soc_videosoc_sdram_bankmachine4_refresh_req) begin
				vns_bankmachine4_next_state <= 2'd3;
			end else begin
				if (soc_videosoc_sdram_bankmachine4_source_valid) begin
					if (soc_videosoc_sdram_bankmachine4_has_openrow) begin
						if (soc_videosoc_sdram_bankmachine4_hit) begin
							soc_videosoc_sdram_bankmachine4_cmd_valid <= 1'd1;
							if (soc_videosoc_sdram_bankmachine4_source_payload_we) begin
								soc_videosoc_sdram_bankmachine4_req_wdata_ready <= soc_videosoc_sdram_bankmachine4_cmd_ready;
								soc_videosoc_sdram_bankmachine4_cmd_payload_is_write <= 1'd1;
								soc_videosoc_sdram_bankmachine4_cmd_payload_we <= 1'd1;
							end else begin
								soc_videosoc_sdram_bankmachine4_req_rdata_valid <= soc_videosoc_sdram_bankmachine4_cmd_ready;
								soc_videosoc_sdram_bankmachine4_cmd_payload_is_read <= 1'd1;
							end
							soc_videosoc_sdram_bankmachine4_cmd_payload_cas <= 1'd1;
						end else begin
							vns_bankmachine4_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine4_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign soc_videosoc_sdram_bankmachine5_sink_valid = soc_videosoc_sdram_bankmachine5_req_valid;
assign soc_videosoc_sdram_bankmachine5_req_ready = soc_videosoc_sdram_bankmachine5_sink_ready;
assign soc_videosoc_sdram_bankmachine5_sink_payload_we = soc_videosoc_sdram_bankmachine5_req_we;
assign soc_videosoc_sdram_bankmachine5_sink_payload_adr = soc_videosoc_sdram_bankmachine5_req_adr;
assign soc_videosoc_sdram_bankmachine5_source_ready = (soc_videosoc_sdram_bankmachine5_req_wdata_ready | soc_videosoc_sdram_bankmachine5_req_rdata_valid);
assign soc_videosoc_sdram_bankmachine5_req_lock = soc_videosoc_sdram_bankmachine5_source_valid;
assign soc_videosoc_sdram_bankmachine5_hit = (soc_videosoc_sdram_bankmachine5_openrow == soc_videosoc_sdram_bankmachine5_source_payload_adr[21:7]);
assign soc_videosoc_sdram_bankmachine5_cmd_payload_ba = 3'd5;
always @(*) begin
	soc_videosoc_sdram_bankmachine5_cmd_payload_a <= 15'd0;
	if (soc_videosoc_sdram_bankmachine5_sel_row_adr) begin
		soc_videosoc_sdram_bankmachine5_cmd_payload_a <= soc_videosoc_sdram_bankmachine5_source_payload_adr[21:7];
	end else begin
		soc_videosoc_sdram_bankmachine5_cmd_payload_a <= {soc_videosoc_sdram_bankmachine5_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign soc_videosoc_sdram_bankmachine5_wait = (~((soc_videosoc_sdram_bankmachine5_cmd_valid & soc_videosoc_sdram_bankmachine5_cmd_ready) & soc_videosoc_sdram_bankmachine5_cmd_payload_is_write));
assign soc_videosoc_sdram_bankmachine5_syncfifo5_din = {soc_videosoc_sdram_bankmachine5_fifo_in_last, soc_videosoc_sdram_bankmachine5_fifo_in_first, soc_videosoc_sdram_bankmachine5_fifo_in_payload_adr, soc_videosoc_sdram_bankmachine5_fifo_in_payload_we};
assign {soc_videosoc_sdram_bankmachine5_fifo_out_last, soc_videosoc_sdram_bankmachine5_fifo_out_first, soc_videosoc_sdram_bankmachine5_fifo_out_payload_adr, soc_videosoc_sdram_bankmachine5_fifo_out_payload_we} = soc_videosoc_sdram_bankmachine5_syncfifo5_dout;
assign soc_videosoc_sdram_bankmachine5_sink_ready = soc_videosoc_sdram_bankmachine5_syncfifo5_writable;
assign soc_videosoc_sdram_bankmachine5_syncfifo5_we = soc_videosoc_sdram_bankmachine5_sink_valid;
assign soc_videosoc_sdram_bankmachine5_fifo_in_first = soc_videosoc_sdram_bankmachine5_sink_first;
assign soc_videosoc_sdram_bankmachine5_fifo_in_last = soc_videosoc_sdram_bankmachine5_sink_last;
assign soc_videosoc_sdram_bankmachine5_fifo_in_payload_we = soc_videosoc_sdram_bankmachine5_sink_payload_we;
assign soc_videosoc_sdram_bankmachine5_fifo_in_payload_adr = soc_videosoc_sdram_bankmachine5_sink_payload_adr;
assign soc_videosoc_sdram_bankmachine5_source_valid = soc_videosoc_sdram_bankmachine5_syncfifo5_readable;
assign soc_videosoc_sdram_bankmachine5_source_first = soc_videosoc_sdram_bankmachine5_fifo_out_first;
assign soc_videosoc_sdram_bankmachine5_source_last = soc_videosoc_sdram_bankmachine5_fifo_out_last;
assign soc_videosoc_sdram_bankmachine5_source_payload_we = soc_videosoc_sdram_bankmachine5_fifo_out_payload_we;
assign soc_videosoc_sdram_bankmachine5_source_payload_adr = soc_videosoc_sdram_bankmachine5_fifo_out_payload_adr;
assign soc_videosoc_sdram_bankmachine5_syncfifo5_re = soc_videosoc_sdram_bankmachine5_source_ready;
always @(*) begin
	soc_videosoc_sdram_bankmachine5_wrport_adr <= 3'd0;
	if (soc_videosoc_sdram_bankmachine5_replace) begin
		soc_videosoc_sdram_bankmachine5_wrport_adr <= (soc_videosoc_sdram_bankmachine5_produce - 1'd1);
	end else begin
		soc_videosoc_sdram_bankmachine5_wrport_adr <= soc_videosoc_sdram_bankmachine5_produce;
	end
end
assign soc_videosoc_sdram_bankmachine5_wrport_dat_w = soc_videosoc_sdram_bankmachine5_syncfifo5_din;
assign soc_videosoc_sdram_bankmachine5_wrport_we = (soc_videosoc_sdram_bankmachine5_syncfifo5_we & (soc_videosoc_sdram_bankmachine5_syncfifo5_writable | soc_videosoc_sdram_bankmachine5_replace));
assign soc_videosoc_sdram_bankmachine5_do_read = (soc_videosoc_sdram_bankmachine5_syncfifo5_readable & soc_videosoc_sdram_bankmachine5_syncfifo5_re);
assign soc_videosoc_sdram_bankmachine5_rdport_adr = soc_videosoc_sdram_bankmachine5_consume;
assign soc_videosoc_sdram_bankmachine5_syncfifo5_dout = soc_videosoc_sdram_bankmachine5_rdport_dat_r;
assign soc_videosoc_sdram_bankmachine5_syncfifo5_writable = (soc_videosoc_sdram_bankmachine5_level != 4'd8);
assign soc_videosoc_sdram_bankmachine5_syncfifo5_readable = (soc_videosoc_sdram_bankmachine5_level != 1'd0);
assign soc_videosoc_sdram_bankmachine5_done = (soc_videosoc_sdram_bankmachine5_count == 1'd0);
always @(*) begin
	soc_videosoc_sdram_bankmachine5_track_open <= 1'd0;
	soc_videosoc_sdram_bankmachine5_track_close <= 1'd0;
	soc_videosoc_sdram_bankmachine5_cmd_payload_cas <= 1'd0;
	soc_videosoc_sdram_bankmachine5_cmd_payload_ras <= 1'd0;
	soc_videosoc_sdram_bankmachine5_cmd_payload_we <= 1'd0;
	soc_videosoc_sdram_bankmachine5_sel_row_adr <= 1'd0;
	soc_videosoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd0;
	soc_videosoc_sdram_bankmachine5_cmd_payload_is_read <= 1'd0;
	soc_videosoc_sdram_bankmachine5_cmd_payload_is_write <= 1'd0;
	soc_videosoc_sdram_bankmachine5_req_wdata_ready <= 1'd0;
	soc_videosoc_sdram_bankmachine5_req_rdata_valid <= 1'd0;
	soc_videosoc_sdram_bankmachine5_refresh_gnt <= 1'd0;
	soc_videosoc_sdram_bankmachine5_cmd_valid <= 1'd0;
	vns_bankmachine5_next_state <= 3'd0;
	vns_bankmachine5_next_state <= vns_bankmachine5_state;
	case (vns_bankmachine5_state)
		1'd1: begin
			if (soc_videosoc_sdram_bankmachine5_done) begin
				soc_videosoc_sdram_bankmachine5_cmd_valid <= 1'd1;
				if (soc_videosoc_sdram_bankmachine5_cmd_ready) begin
					vns_bankmachine5_next_state <= 3'd4;
				end
				soc_videosoc_sdram_bankmachine5_cmd_payload_ras <= 1'd1;
				soc_videosoc_sdram_bankmachine5_cmd_payload_we <= 1'd1;
				soc_videosoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine5_track_close <= 1'd1;
		end
		2'd2: begin
			soc_videosoc_sdram_bankmachine5_sel_row_adr <= 1'd1;
			soc_videosoc_sdram_bankmachine5_track_open <= 1'd1;
			soc_videosoc_sdram_bankmachine5_cmd_valid <= 1'd1;
			soc_videosoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd1;
			if (soc_videosoc_sdram_bankmachine5_cmd_ready) begin
				vns_bankmachine5_next_state <= 3'd6;
			end
			soc_videosoc_sdram_bankmachine5_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (soc_videosoc_sdram_bankmachine5_done) begin
				soc_videosoc_sdram_bankmachine5_refresh_gnt <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine5_track_close <= 1'd1;
			soc_videosoc_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videosoc_sdram_bankmachine5_refresh_req)) begin
				vns_bankmachine5_next_state <= 1'd0;
			end
		end
		3'd4: begin
			vns_bankmachine5_next_state <= 3'd5;
		end
		3'd5: begin
			vns_bankmachine5_next_state <= 2'd2;
		end
		3'd6: begin
			vns_bankmachine5_next_state <= 3'd7;
		end
		3'd7: begin
			vns_bankmachine5_next_state <= 1'd0;
		end
		default: begin
			if (soc_videosoc_sdram_bankmachine5_refresh_req) begin
				vns_bankmachine5_next_state <= 2'd3;
			end else begin
				if (soc_videosoc_sdram_bankmachine5_source_valid) begin
					if (soc_videosoc_sdram_bankmachine5_has_openrow) begin
						if (soc_videosoc_sdram_bankmachine5_hit) begin
							soc_videosoc_sdram_bankmachine5_cmd_valid <= 1'd1;
							if (soc_videosoc_sdram_bankmachine5_source_payload_we) begin
								soc_videosoc_sdram_bankmachine5_req_wdata_ready <= soc_videosoc_sdram_bankmachine5_cmd_ready;
								soc_videosoc_sdram_bankmachine5_cmd_payload_is_write <= 1'd1;
								soc_videosoc_sdram_bankmachine5_cmd_payload_we <= 1'd1;
							end else begin
								soc_videosoc_sdram_bankmachine5_req_rdata_valid <= soc_videosoc_sdram_bankmachine5_cmd_ready;
								soc_videosoc_sdram_bankmachine5_cmd_payload_is_read <= 1'd1;
							end
							soc_videosoc_sdram_bankmachine5_cmd_payload_cas <= 1'd1;
						end else begin
							vns_bankmachine5_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine5_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign soc_videosoc_sdram_bankmachine6_sink_valid = soc_videosoc_sdram_bankmachine6_req_valid;
assign soc_videosoc_sdram_bankmachine6_req_ready = soc_videosoc_sdram_bankmachine6_sink_ready;
assign soc_videosoc_sdram_bankmachine6_sink_payload_we = soc_videosoc_sdram_bankmachine6_req_we;
assign soc_videosoc_sdram_bankmachine6_sink_payload_adr = soc_videosoc_sdram_bankmachine6_req_adr;
assign soc_videosoc_sdram_bankmachine6_source_ready = (soc_videosoc_sdram_bankmachine6_req_wdata_ready | soc_videosoc_sdram_bankmachine6_req_rdata_valid);
assign soc_videosoc_sdram_bankmachine6_req_lock = soc_videosoc_sdram_bankmachine6_source_valid;
assign soc_videosoc_sdram_bankmachine6_hit = (soc_videosoc_sdram_bankmachine6_openrow == soc_videosoc_sdram_bankmachine6_source_payload_adr[21:7]);
assign soc_videosoc_sdram_bankmachine6_cmd_payload_ba = 3'd6;
always @(*) begin
	soc_videosoc_sdram_bankmachine6_cmd_payload_a <= 15'd0;
	if (soc_videosoc_sdram_bankmachine6_sel_row_adr) begin
		soc_videosoc_sdram_bankmachine6_cmd_payload_a <= soc_videosoc_sdram_bankmachine6_source_payload_adr[21:7];
	end else begin
		soc_videosoc_sdram_bankmachine6_cmd_payload_a <= {soc_videosoc_sdram_bankmachine6_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign soc_videosoc_sdram_bankmachine6_wait = (~((soc_videosoc_sdram_bankmachine6_cmd_valid & soc_videosoc_sdram_bankmachine6_cmd_ready) & soc_videosoc_sdram_bankmachine6_cmd_payload_is_write));
assign soc_videosoc_sdram_bankmachine6_syncfifo6_din = {soc_videosoc_sdram_bankmachine6_fifo_in_last, soc_videosoc_sdram_bankmachine6_fifo_in_first, soc_videosoc_sdram_bankmachine6_fifo_in_payload_adr, soc_videosoc_sdram_bankmachine6_fifo_in_payload_we};
assign {soc_videosoc_sdram_bankmachine6_fifo_out_last, soc_videosoc_sdram_bankmachine6_fifo_out_first, soc_videosoc_sdram_bankmachine6_fifo_out_payload_adr, soc_videosoc_sdram_bankmachine6_fifo_out_payload_we} = soc_videosoc_sdram_bankmachine6_syncfifo6_dout;
assign soc_videosoc_sdram_bankmachine6_sink_ready = soc_videosoc_sdram_bankmachine6_syncfifo6_writable;
assign soc_videosoc_sdram_bankmachine6_syncfifo6_we = soc_videosoc_sdram_bankmachine6_sink_valid;
assign soc_videosoc_sdram_bankmachine6_fifo_in_first = soc_videosoc_sdram_bankmachine6_sink_first;
assign soc_videosoc_sdram_bankmachine6_fifo_in_last = soc_videosoc_sdram_bankmachine6_sink_last;
assign soc_videosoc_sdram_bankmachine6_fifo_in_payload_we = soc_videosoc_sdram_bankmachine6_sink_payload_we;
assign soc_videosoc_sdram_bankmachine6_fifo_in_payload_adr = soc_videosoc_sdram_bankmachine6_sink_payload_adr;
assign soc_videosoc_sdram_bankmachine6_source_valid = soc_videosoc_sdram_bankmachine6_syncfifo6_readable;
assign soc_videosoc_sdram_bankmachine6_source_first = soc_videosoc_sdram_bankmachine6_fifo_out_first;
assign soc_videosoc_sdram_bankmachine6_source_last = soc_videosoc_sdram_bankmachine6_fifo_out_last;
assign soc_videosoc_sdram_bankmachine6_source_payload_we = soc_videosoc_sdram_bankmachine6_fifo_out_payload_we;
assign soc_videosoc_sdram_bankmachine6_source_payload_adr = soc_videosoc_sdram_bankmachine6_fifo_out_payload_adr;
assign soc_videosoc_sdram_bankmachine6_syncfifo6_re = soc_videosoc_sdram_bankmachine6_source_ready;
always @(*) begin
	soc_videosoc_sdram_bankmachine6_wrport_adr <= 3'd0;
	if (soc_videosoc_sdram_bankmachine6_replace) begin
		soc_videosoc_sdram_bankmachine6_wrport_adr <= (soc_videosoc_sdram_bankmachine6_produce - 1'd1);
	end else begin
		soc_videosoc_sdram_bankmachine6_wrport_adr <= soc_videosoc_sdram_bankmachine6_produce;
	end
end
assign soc_videosoc_sdram_bankmachine6_wrport_dat_w = soc_videosoc_sdram_bankmachine6_syncfifo6_din;
assign soc_videosoc_sdram_bankmachine6_wrport_we = (soc_videosoc_sdram_bankmachine6_syncfifo6_we & (soc_videosoc_sdram_bankmachine6_syncfifo6_writable | soc_videosoc_sdram_bankmachine6_replace));
assign soc_videosoc_sdram_bankmachine6_do_read = (soc_videosoc_sdram_bankmachine6_syncfifo6_readable & soc_videosoc_sdram_bankmachine6_syncfifo6_re);
assign soc_videosoc_sdram_bankmachine6_rdport_adr = soc_videosoc_sdram_bankmachine6_consume;
assign soc_videosoc_sdram_bankmachine6_syncfifo6_dout = soc_videosoc_sdram_bankmachine6_rdport_dat_r;
assign soc_videosoc_sdram_bankmachine6_syncfifo6_writable = (soc_videosoc_sdram_bankmachine6_level != 4'd8);
assign soc_videosoc_sdram_bankmachine6_syncfifo6_readable = (soc_videosoc_sdram_bankmachine6_level != 1'd0);
assign soc_videosoc_sdram_bankmachine6_done = (soc_videosoc_sdram_bankmachine6_count == 1'd0);
always @(*) begin
	soc_videosoc_sdram_bankmachine6_refresh_gnt <= 1'd0;
	soc_videosoc_sdram_bankmachine6_cmd_valid <= 1'd0;
	soc_videosoc_sdram_bankmachine6_track_open <= 1'd0;
	soc_videosoc_sdram_bankmachine6_track_close <= 1'd0;
	soc_videosoc_sdram_bankmachine6_cmd_payload_cas <= 1'd0;
	soc_videosoc_sdram_bankmachine6_cmd_payload_ras <= 1'd0;
	vns_bankmachine6_next_state <= 3'd0;
	soc_videosoc_sdram_bankmachine6_cmd_payload_we <= 1'd0;
	soc_videosoc_sdram_bankmachine6_sel_row_adr <= 1'd0;
	soc_videosoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd0;
	soc_videosoc_sdram_bankmachine6_cmd_payload_is_read <= 1'd0;
	soc_videosoc_sdram_bankmachine6_cmd_payload_is_write <= 1'd0;
	soc_videosoc_sdram_bankmachine6_req_wdata_ready <= 1'd0;
	soc_videosoc_sdram_bankmachine6_req_rdata_valid <= 1'd0;
	vns_bankmachine6_next_state <= vns_bankmachine6_state;
	case (vns_bankmachine6_state)
		1'd1: begin
			if (soc_videosoc_sdram_bankmachine6_done) begin
				soc_videosoc_sdram_bankmachine6_cmd_valid <= 1'd1;
				if (soc_videosoc_sdram_bankmachine6_cmd_ready) begin
					vns_bankmachine6_next_state <= 3'd4;
				end
				soc_videosoc_sdram_bankmachine6_cmd_payload_ras <= 1'd1;
				soc_videosoc_sdram_bankmachine6_cmd_payload_we <= 1'd1;
				soc_videosoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine6_track_close <= 1'd1;
		end
		2'd2: begin
			soc_videosoc_sdram_bankmachine6_sel_row_adr <= 1'd1;
			soc_videosoc_sdram_bankmachine6_track_open <= 1'd1;
			soc_videosoc_sdram_bankmachine6_cmd_valid <= 1'd1;
			soc_videosoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd1;
			if (soc_videosoc_sdram_bankmachine6_cmd_ready) begin
				vns_bankmachine6_next_state <= 3'd6;
			end
			soc_videosoc_sdram_bankmachine6_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (soc_videosoc_sdram_bankmachine6_done) begin
				soc_videosoc_sdram_bankmachine6_refresh_gnt <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine6_track_close <= 1'd1;
			soc_videosoc_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videosoc_sdram_bankmachine6_refresh_req)) begin
				vns_bankmachine6_next_state <= 1'd0;
			end
		end
		3'd4: begin
			vns_bankmachine6_next_state <= 3'd5;
		end
		3'd5: begin
			vns_bankmachine6_next_state <= 2'd2;
		end
		3'd6: begin
			vns_bankmachine6_next_state <= 3'd7;
		end
		3'd7: begin
			vns_bankmachine6_next_state <= 1'd0;
		end
		default: begin
			if (soc_videosoc_sdram_bankmachine6_refresh_req) begin
				vns_bankmachine6_next_state <= 2'd3;
			end else begin
				if (soc_videosoc_sdram_bankmachine6_source_valid) begin
					if (soc_videosoc_sdram_bankmachine6_has_openrow) begin
						if (soc_videosoc_sdram_bankmachine6_hit) begin
							soc_videosoc_sdram_bankmachine6_cmd_valid <= 1'd1;
							if (soc_videosoc_sdram_bankmachine6_source_payload_we) begin
								soc_videosoc_sdram_bankmachine6_req_wdata_ready <= soc_videosoc_sdram_bankmachine6_cmd_ready;
								soc_videosoc_sdram_bankmachine6_cmd_payload_is_write <= 1'd1;
								soc_videosoc_sdram_bankmachine6_cmd_payload_we <= 1'd1;
							end else begin
								soc_videosoc_sdram_bankmachine6_req_rdata_valid <= soc_videosoc_sdram_bankmachine6_cmd_ready;
								soc_videosoc_sdram_bankmachine6_cmd_payload_is_read <= 1'd1;
							end
							soc_videosoc_sdram_bankmachine6_cmd_payload_cas <= 1'd1;
						end else begin
							vns_bankmachine6_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine6_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign soc_videosoc_sdram_bankmachine7_sink_valid = soc_videosoc_sdram_bankmachine7_req_valid;
assign soc_videosoc_sdram_bankmachine7_req_ready = soc_videosoc_sdram_bankmachine7_sink_ready;
assign soc_videosoc_sdram_bankmachine7_sink_payload_we = soc_videosoc_sdram_bankmachine7_req_we;
assign soc_videosoc_sdram_bankmachine7_sink_payload_adr = soc_videosoc_sdram_bankmachine7_req_adr;
assign soc_videosoc_sdram_bankmachine7_source_ready = (soc_videosoc_sdram_bankmachine7_req_wdata_ready | soc_videosoc_sdram_bankmachine7_req_rdata_valid);
assign soc_videosoc_sdram_bankmachine7_req_lock = soc_videosoc_sdram_bankmachine7_source_valid;
assign soc_videosoc_sdram_bankmachine7_hit = (soc_videosoc_sdram_bankmachine7_openrow == soc_videosoc_sdram_bankmachine7_source_payload_adr[21:7]);
assign soc_videosoc_sdram_bankmachine7_cmd_payload_ba = 3'd7;
always @(*) begin
	soc_videosoc_sdram_bankmachine7_cmd_payload_a <= 15'd0;
	if (soc_videosoc_sdram_bankmachine7_sel_row_adr) begin
		soc_videosoc_sdram_bankmachine7_cmd_payload_a <= soc_videosoc_sdram_bankmachine7_source_payload_adr[21:7];
	end else begin
		soc_videosoc_sdram_bankmachine7_cmd_payload_a <= {soc_videosoc_sdram_bankmachine7_source_payload_adr[6:0], {3{1'd0}}};
	end
end
assign soc_videosoc_sdram_bankmachine7_wait = (~((soc_videosoc_sdram_bankmachine7_cmd_valid & soc_videosoc_sdram_bankmachine7_cmd_ready) & soc_videosoc_sdram_bankmachine7_cmd_payload_is_write));
assign soc_videosoc_sdram_bankmachine7_syncfifo7_din = {soc_videosoc_sdram_bankmachine7_fifo_in_last, soc_videosoc_sdram_bankmachine7_fifo_in_first, soc_videosoc_sdram_bankmachine7_fifo_in_payload_adr, soc_videosoc_sdram_bankmachine7_fifo_in_payload_we};
assign {soc_videosoc_sdram_bankmachine7_fifo_out_last, soc_videosoc_sdram_bankmachine7_fifo_out_first, soc_videosoc_sdram_bankmachine7_fifo_out_payload_adr, soc_videosoc_sdram_bankmachine7_fifo_out_payload_we} = soc_videosoc_sdram_bankmachine7_syncfifo7_dout;
assign soc_videosoc_sdram_bankmachine7_sink_ready = soc_videosoc_sdram_bankmachine7_syncfifo7_writable;
assign soc_videosoc_sdram_bankmachine7_syncfifo7_we = soc_videosoc_sdram_bankmachine7_sink_valid;
assign soc_videosoc_sdram_bankmachine7_fifo_in_first = soc_videosoc_sdram_bankmachine7_sink_first;
assign soc_videosoc_sdram_bankmachine7_fifo_in_last = soc_videosoc_sdram_bankmachine7_sink_last;
assign soc_videosoc_sdram_bankmachine7_fifo_in_payload_we = soc_videosoc_sdram_bankmachine7_sink_payload_we;
assign soc_videosoc_sdram_bankmachine7_fifo_in_payload_adr = soc_videosoc_sdram_bankmachine7_sink_payload_adr;
assign soc_videosoc_sdram_bankmachine7_source_valid = soc_videosoc_sdram_bankmachine7_syncfifo7_readable;
assign soc_videosoc_sdram_bankmachine7_source_first = soc_videosoc_sdram_bankmachine7_fifo_out_first;
assign soc_videosoc_sdram_bankmachine7_source_last = soc_videosoc_sdram_bankmachine7_fifo_out_last;
assign soc_videosoc_sdram_bankmachine7_source_payload_we = soc_videosoc_sdram_bankmachine7_fifo_out_payload_we;
assign soc_videosoc_sdram_bankmachine7_source_payload_adr = soc_videosoc_sdram_bankmachine7_fifo_out_payload_adr;
assign soc_videosoc_sdram_bankmachine7_syncfifo7_re = soc_videosoc_sdram_bankmachine7_source_ready;
always @(*) begin
	soc_videosoc_sdram_bankmachine7_wrport_adr <= 3'd0;
	if (soc_videosoc_sdram_bankmachine7_replace) begin
		soc_videosoc_sdram_bankmachine7_wrport_adr <= (soc_videosoc_sdram_bankmachine7_produce - 1'd1);
	end else begin
		soc_videosoc_sdram_bankmachine7_wrport_adr <= soc_videosoc_sdram_bankmachine7_produce;
	end
end
assign soc_videosoc_sdram_bankmachine7_wrport_dat_w = soc_videosoc_sdram_bankmachine7_syncfifo7_din;
assign soc_videosoc_sdram_bankmachine7_wrport_we = (soc_videosoc_sdram_bankmachine7_syncfifo7_we & (soc_videosoc_sdram_bankmachine7_syncfifo7_writable | soc_videosoc_sdram_bankmachine7_replace));
assign soc_videosoc_sdram_bankmachine7_do_read = (soc_videosoc_sdram_bankmachine7_syncfifo7_readable & soc_videosoc_sdram_bankmachine7_syncfifo7_re);
assign soc_videosoc_sdram_bankmachine7_rdport_adr = soc_videosoc_sdram_bankmachine7_consume;
assign soc_videosoc_sdram_bankmachine7_syncfifo7_dout = soc_videosoc_sdram_bankmachine7_rdport_dat_r;
assign soc_videosoc_sdram_bankmachine7_syncfifo7_writable = (soc_videosoc_sdram_bankmachine7_level != 4'd8);
assign soc_videosoc_sdram_bankmachine7_syncfifo7_readable = (soc_videosoc_sdram_bankmachine7_level != 1'd0);
assign soc_videosoc_sdram_bankmachine7_done = (soc_videosoc_sdram_bankmachine7_count == 1'd0);
always @(*) begin
	soc_videosoc_sdram_bankmachine7_cmd_payload_we <= 1'd0;
	soc_videosoc_sdram_bankmachine7_sel_row_adr <= 1'd0;
	soc_videosoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd0;
	soc_videosoc_sdram_bankmachine7_cmd_payload_is_read <= 1'd0;
	soc_videosoc_sdram_bankmachine7_cmd_payload_is_write <= 1'd0;
	soc_videosoc_sdram_bankmachine7_req_wdata_ready <= 1'd0;
	soc_videosoc_sdram_bankmachine7_req_rdata_valid <= 1'd0;
	soc_videosoc_sdram_bankmachine7_refresh_gnt <= 1'd0;
	soc_videosoc_sdram_bankmachine7_cmd_valid <= 1'd0;
	vns_bankmachine7_next_state <= 3'd0;
	soc_videosoc_sdram_bankmachine7_cmd_payload_cas <= 1'd0;
	soc_videosoc_sdram_bankmachine7_track_open <= 1'd0;
	soc_videosoc_sdram_bankmachine7_track_close <= 1'd0;
	soc_videosoc_sdram_bankmachine7_cmd_payload_ras <= 1'd0;
	vns_bankmachine7_next_state <= vns_bankmachine7_state;
	case (vns_bankmachine7_state)
		1'd1: begin
			if (soc_videosoc_sdram_bankmachine7_done) begin
				soc_videosoc_sdram_bankmachine7_cmd_valid <= 1'd1;
				if (soc_videosoc_sdram_bankmachine7_cmd_ready) begin
					vns_bankmachine7_next_state <= 3'd4;
				end
				soc_videosoc_sdram_bankmachine7_cmd_payload_ras <= 1'd1;
				soc_videosoc_sdram_bankmachine7_cmd_payload_we <= 1'd1;
				soc_videosoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine7_track_close <= 1'd1;
		end
		2'd2: begin
			soc_videosoc_sdram_bankmachine7_sel_row_adr <= 1'd1;
			soc_videosoc_sdram_bankmachine7_track_open <= 1'd1;
			soc_videosoc_sdram_bankmachine7_cmd_valid <= 1'd1;
			soc_videosoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd1;
			if (soc_videosoc_sdram_bankmachine7_cmd_ready) begin
				vns_bankmachine7_next_state <= 3'd6;
			end
			soc_videosoc_sdram_bankmachine7_cmd_payload_ras <= 1'd1;
		end
		2'd3: begin
			if (soc_videosoc_sdram_bankmachine7_done) begin
				soc_videosoc_sdram_bankmachine7_refresh_gnt <= 1'd1;
			end
			soc_videosoc_sdram_bankmachine7_track_close <= 1'd1;
			soc_videosoc_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd1;
			if ((~soc_videosoc_sdram_bankmachine7_refresh_req)) begin
				vns_bankmachine7_next_state <= 1'd0;
			end
		end
		3'd4: begin
			vns_bankmachine7_next_state <= 3'd5;
		end
		3'd5: begin
			vns_bankmachine7_next_state <= 2'd2;
		end
		3'd6: begin
			vns_bankmachine7_next_state <= 3'd7;
		end
		3'd7: begin
			vns_bankmachine7_next_state <= 1'd0;
		end
		default: begin
			if (soc_videosoc_sdram_bankmachine7_refresh_req) begin
				vns_bankmachine7_next_state <= 2'd3;
			end else begin
				if (soc_videosoc_sdram_bankmachine7_source_valid) begin
					if (soc_videosoc_sdram_bankmachine7_has_openrow) begin
						if (soc_videosoc_sdram_bankmachine7_hit) begin
							soc_videosoc_sdram_bankmachine7_cmd_valid <= 1'd1;
							if (soc_videosoc_sdram_bankmachine7_source_payload_we) begin
								soc_videosoc_sdram_bankmachine7_req_wdata_ready <= soc_videosoc_sdram_bankmachine7_cmd_ready;
								soc_videosoc_sdram_bankmachine7_cmd_payload_is_write <= 1'd1;
								soc_videosoc_sdram_bankmachine7_cmd_payload_we <= 1'd1;
							end else begin
								soc_videosoc_sdram_bankmachine7_req_rdata_valid <= soc_videosoc_sdram_bankmachine7_cmd_ready;
								soc_videosoc_sdram_bankmachine7_cmd_payload_is_read <= 1'd1;
							end
							soc_videosoc_sdram_bankmachine7_cmd_payload_cas <= 1'd1;
						end else begin
							vns_bankmachine7_next_state <= 1'd1;
						end
					end else begin
						vns_bankmachine7_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign soc_videosoc_sdram_read_available = ((((((((soc_videosoc_sdram_bankmachine0_cmd_valid & soc_videosoc_sdram_bankmachine0_cmd_payload_is_read) | (soc_videosoc_sdram_bankmachine1_cmd_valid & soc_videosoc_sdram_bankmachine1_cmd_payload_is_read)) | (soc_videosoc_sdram_bankmachine2_cmd_valid & soc_videosoc_sdram_bankmachine2_cmd_payload_is_read)) | (soc_videosoc_sdram_bankmachine3_cmd_valid & soc_videosoc_sdram_bankmachine3_cmd_payload_is_read)) | (soc_videosoc_sdram_bankmachine4_cmd_valid & soc_videosoc_sdram_bankmachine4_cmd_payload_is_read)) | (soc_videosoc_sdram_bankmachine5_cmd_valid & soc_videosoc_sdram_bankmachine5_cmd_payload_is_read)) | (soc_videosoc_sdram_bankmachine6_cmd_valid & soc_videosoc_sdram_bankmachine6_cmd_payload_is_read)) | (soc_videosoc_sdram_bankmachine7_cmd_valid & soc_videosoc_sdram_bankmachine7_cmd_payload_is_read));
assign soc_videosoc_sdram_write_available = ((((((((soc_videosoc_sdram_bankmachine0_cmd_valid & soc_videosoc_sdram_bankmachine0_cmd_payload_is_write) | (soc_videosoc_sdram_bankmachine1_cmd_valid & soc_videosoc_sdram_bankmachine1_cmd_payload_is_write)) | (soc_videosoc_sdram_bankmachine2_cmd_valid & soc_videosoc_sdram_bankmachine2_cmd_payload_is_write)) | (soc_videosoc_sdram_bankmachine3_cmd_valid & soc_videosoc_sdram_bankmachine3_cmd_payload_is_write)) | (soc_videosoc_sdram_bankmachine4_cmd_valid & soc_videosoc_sdram_bankmachine4_cmd_payload_is_write)) | (soc_videosoc_sdram_bankmachine5_cmd_valid & soc_videosoc_sdram_bankmachine5_cmd_payload_is_write)) | (soc_videosoc_sdram_bankmachine6_cmd_valid & soc_videosoc_sdram_bankmachine6_cmd_payload_is_write)) | (soc_videosoc_sdram_bankmachine7_cmd_valid & soc_videosoc_sdram_bankmachine7_cmd_payload_is_write));
assign soc_videosoc_sdram_max_time0 = (soc_videosoc_sdram_time0 == 1'd0);
assign soc_videosoc_sdram_max_time1 = (soc_videosoc_sdram_time1 == 1'd0);
assign soc_videosoc_sdram_bankmachine0_refresh_req = soc_videosoc_sdram_cmd_valid;
assign soc_videosoc_sdram_bankmachine1_refresh_req = soc_videosoc_sdram_cmd_valid;
assign soc_videosoc_sdram_bankmachine2_refresh_req = soc_videosoc_sdram_cmd_valid;
assign soc_videosoc_sdram_bankmachine3_refresh_req = soc_videosoc_sdram_cmd_valid;
assign soc_videosoc_sdram_bankmachine4_refresh_req = soc_videosoc_sdram_cmd_valid;
assign soc_videosoc_sdram_bankmachine5_refresh_req = soc_videosoc_sdram_cmd_valid;
assign soc_videosoc_sdram_bankmachine6_refresh_req = soc_videosoc_sdram_cmd_valid;
assign soc_videosoc_sdram_bankmachine7_refresh_req = soc_videosoc_sdram_cmd_valid;
assign soc_videosoc_sdram_go_to_refresh = (((((((soc_videosoc_sdram_bankmachine0_refresh_gnt & soc_videosoc_sdram_bankmachine1_refresh_gnt) & soc_videosoc_sdram_bankmachine2_refresh_gnt) & soc_videosoc_sdram_bankmachine3_refresh_gnt) & soc_videosoc_sdram_bankmachine4_refresh_gnt) & soc_videosoc_sdram_bankmachine5_refresh_gnt) & soc_videosoc_sdram_bankmachine6_refresh_gnt) & soc_videosoc_sdram_bankmachine7_refresh_gnt);
assign soc_videosoc_sdram_interface_rdata = {soc_videosoc_sdram_dfi_p3_rddata, soc_videosoc_sdram_dfi_p2_rddata, soc_videosoc_sdram_dfi_p1_rddata, soc_videosoc_sdram_dfi_p0_rddata};
assign {soc_videosoc_sdram_dfi_p3_wrdata, soc_videosoc_sdram_dfi_p2_wrdata, soc_videosoc_sdram_dfi_p1_wrdata, soc_videosoc_sdram_dfi_p0_wrdata} = soc_videosoc_sdram_interface_wdata;
assign {soc_videosoc_sdram_dfi_p3_wrdata_mask, soc_videosoc_sdram_dfi_p2_wrdata_mask, soc_videosoc_sdram_dfi_p1_wrdata_mask, soc_videosoc_sdram_dfi_p0_wrdata_mask} = (~soc_videosoc_sdram_interface_wdata_we);
always @(*) begin
	soc_videosoc_sdram_choose_cmd_valids <= 8'd0;
	soc_videosoc_sdram_choose_cmd_valids[0] <= (soc_videosoc_sdram_bankmachine0_cmd_valid & ((soc_videosoc_sdram_bankmachine0_cmd_payload_is_cmd & soc_videosoc_sdram_choose_cmd_want_cmds) | ((soc_videosoc_sdram_bankmachine0_cmd_payload_is_read == soc_videosoc_sdram_choose_cmd_want_reads) & (soc_videosoc_sdram_bankmachine0_cmd_payload_is_write == soc_videosoc_sdram_choose_cmd_want_writes))));
	soc_videosoc_sdram_choose_cmd_valids[1] <= (soc_videosoc_sdram_bankmachine1_cmd_valid & ((soc_videosoc_sdram_bankmachine1_cmd_payload_is_cmd & soc_videosoc_sdram_choose_cmd_want_cmds) | ((soc_videosoc_sdram_bankmachine1_cmd_payload_is_read == soc_videosoc_sdram_choose_cmd_want_reads) & (soc_videosoc_sdram_bankmachine1_cmd_payload_is_write == soc_videosoc_sdram_choose_cmd_want_writes))));
	soc_videosoc_sdram_choose_cmd_valids[2] <= (soc_videosoc_sdram_bankmachine2_cmd_valid & ((soc_videosoc_sdram_bankmachine2_cmd_payload_is_cmd & soc_videosoc_sdram_choose_cmd_want_cmds) | ((soc_videosoc_sdram_bankmachine2_cmd_payload_is_read == soc_videosoc_sdram_choose_cmd_want_reads) & (soc_videosoc_sdram_bankmachine2_cmd_payload_is_write == soc_videosoc_sdram_choose_cmd_want_writes))));
	soc_videosoc_sdram_choose_cmd_valids[3] <= (soc_videosoc_sdram_bankmachine3_cmd_valid & ((soc_videosoc_sdram_bankmachine3_cmd_payload_is_cmd & soc_videosoc_sdram_choose_cmd_want_cmds) | ((soc_videosoc_sdram_bankmachine3_cmd_payload_is_read == soc_videosoc_sdram_choose_cmd_want_reads) & (soc_videosoc_sdram_bankmachine3_cmd_payload_is_write == soc_videosoc_sdram_choose_cmd_want_writes))));
	soc_videosoc_sdram_choose_cmd_valids[4] <= (soc_videosoc_sdram_bankmachine4_cmd_valid & ((soc_videosoc_sdram_bankmachine4_cmd_payload_is_cmd & soc_videosoc_sdram_choose_cmd_want_cmds) | ((soc_videosoc_sdram_bankmachine4_cmd_payload_is_read == soc_videosoc_sdram_choose_cmd_want_reads) & (soc_videosoc_sdram_bankmachine4_cmd_payload_is_write == soc_videosoc_sdram_choose_cmd_want_writes))));
	soc_videosoc_sdram_choose_cmd_valids[5] <= (soc_videosoc_sdram_bankmachine5_cmd_valid & ((soc_videosoc_sdram_bankmachine5_cmd_payload_is_cmd & soc_videosoc_sdram_choose_cmd_want_cmds) | ((soc_videosoc_sdram_bankmachine5_cmd_payload_is_read == soc_videosoc_sdram_choose_cmd_want_reads) & (soc_videosoc_sdram_bankmachine5_cmd_payload_is_write == soc_videosoc_sdram_choose_cmd_want_writes))));
	soc_videosoc_sdram_choose_cmd_valids[6] <= (soc_videosoc_sdram_bankmachine6_cmd_valid & ((soc_videosoc_sdram_bankmachine6_cmd_payload_is_cmd & soc_videosoc_sdram_choose_cmd_want_cmds) | ((soc_videosoc_sdram_bankmachine6_cmd_payload_is_read == soc_videosoc_sdram_choose_cmd_want_reads) & (soc_videosoc_sdram_bankmachine6_cmd_payload_is_write == soc_videosoc_sdram_choose_cmd_want_writes))));
	soc_videosoc_sdram_choose_cmd_valids[7] <= (soc_videosoc_sdram_bankmachine7_cmd_valid & ((soc_videosoc_sdram_bankmachine7_cmd_payload_is_cmd & soc_videosoc_sdram_choose_cmd_want_cmds) | ((soc_videosoc_sdram_bankmachine7_cmd_payload_is_read == soc_videosoc_sdram_choose_cmd_want_reads) & (soc_videosoc_sdram_bankmachine7_cmd_payload_is_write == soc_videosoc_sdram_choose_cmd_want_writes))));
end
assign soc_videosoc_sdram_choose_cmd_request = soc_videosoc_sdram_choose_cmd_valids;
assign soc_videosoc_sdram_choose_cmd_cmd_valid = vns_comb_rhs_array_muxed0;
assign soc_videosoc_sdram_choose_cmd_cmd_payload_a = vns_comb_rhs_array_muxed1;
assign soc_videosoc_sdram_choose_cmd_cmd_payload_ba = vns_comb_rhs_array_muxed2;
assign soc_videosoc_sdram_choose_cmd_cmd_payload_is_read = vns_comb_rhs_array_muxed3;
assign soc_videosoc_sdram_choose_cmd_cmd_payload_is_write = vns_comb_rhs_array_muxed4;
assign soc_videosoc_sdram_choose_cmd_cmd_payload_is_cmd = vns_comb_rhs_array_muxed5;
always @(*) begin
	soc_videosoc_sdram_choose_cmd_cmd_payload_cas <= 1'd0;
	if (soc_videosoc_sdram_choose_cmd_cmd_valid) begin
		soc_videosoc_sdram_choose_cmd_cmd_payload_cas <= vns_comb_t_array_muxed0;
	end
end
always @(*) begin
	soc_videosoc_sdram_choose_cmd_cmd_payload_ras <= 1'd0;
	if (soc_videosoc_sdram_choose_cmd_cmd_valid) begin
		soc_videosoc_sdram_choose_cmd_cmd_payload_ras <= vns_comb_t_array_muxed1;
	end
end
always @(*) begin
	soc_videosoc_sdram_choose_cmd_cmd_payload_we <= 1'd0;
	if (soc_videosoc_sdram_choose_cmd_cmd_valid) begin
		soc_videosoc_sdram_choose_cmd_cmd_payload_we <= vns_comb_t_array_muxed2;
	end
end
assign soc_videosoc_sdram_choose_cmd_ce = soc_videosoc_sdram_choose_cmd_cmd_ready;
always @(*) begin
	soc_videosoc_sdram_choose_req_valids <= 8'd0;
	soc_videosoc_sdram_choose_req_valids[0] <= (soc_videosoc_sdram_bankmachine0_cmd_valid & ((soc_videosoc_sdram_bankmachine0_cmd_payload_is_cmd & soc_videosoc_sdram_choose_req_want_cmds) | ((soc_videosoc_sdram_bankmachine0_cmd_payload_is_read == soc_videosoc_sdram_choose_req_want_reads) & (soc_videosoc_sdram_bankmachine0_cmd_payload_is_write == soc_videosoc_sdram_choose_req_want_writes))));
	soc_videosoc_sdram_choose_req_valids[1] <= (soc_videosoc_sdram_bankmachine1_cmd_valid & ((soc_videosoc_sdram_bankmachine1_cmd_payload_is_cmd & soc_videosoc_sdram_choose_req_want_cmds) | ((soc_videosoc_sdram_bankmachine1_cmd_payload_is_read == soc_videosoc_sdram_choose_req_want_reads) & (soc_videosoc_sdram_bankmachine1_cmd_payload_is_write == soc_videosoc_sdram_choose_req_want_writes))));
	soc_videosoc_sdram_choose_req_valids[2] <= (soc_videosoc_sdram_bankmachine2_cmd_valid & ((soc_videosoc_sdram_bankmachine2_cmd_payload_is_cmd & soc_videosoc_sdram_choose_req_want_cmds) | ((soc_videosoc_sdram_bankmachine2_cmd_payload_is_read == soc_videosoc_sdram_choose_req_want_reads) & (soc_videosoc_sdram_bankmachine2_cmd_payload_is_write == soc_videosoc_sdram_choose_req_want_writes))));
	soc_videosoc_sdram_choose_req_valids[3] <= (soc_videosoc_sdram_bankmachine3_cmd_valid & ((soc_videosoc_sdram_bankmachine3_cmd_payload_is_cmd & soc_videosoc_sdram_choose_req_want_cmds) | ((soc_videosoc_sdram_bankmachine3_cmd_payload_is_read == soc_videosoc_sdram_choose_req_want_reads) & (soc_videosoc_sdram_bankmachine3_cmd_payload_is_write == soc_videosoc_sdram_choose_req_want_writes))));
	soc_videosoc_sdram_choose_req_valids[4] <= (soc_videosoc_sdram_bankmachine4_cmd_valid & ((soc_videosoc_sdram_bankmachine4_cmd_payload_is_cmd & soc_videosoc_sdram_choose_req_want_cmds) | ((soc_videosoc_sdram_bankmachine4_cmd_payload_is_read == soc_videosoc_sdram_choose_req_want_reads) & (soc_videosoc_sdram_bankmachine4_cmd_payload_is_write == soc_videosoc_sdram_choose_req_want_writes))));
	soc_videosoc_sdram_choose_req_valids[5] <= (soc_videosoc_sdram_bankmachine5_cmd_valid & ((soc_videosoc_sdram_bankmachine5_cmd_payload_is_cmd & soc_videosoc_sdram_choose_req_want_cmds) | ((soc_videosoc_sdram_bankmachine5_cmd_payload_is_read == soc_videosoc_sdram_choose_req_want_reads) & (soc_videosoc_sdram_bankmachine5_cmd_payload_is_write == soc_videosoc_sdram_choose_req_want_writes))));
	soc_videosoc_sdram_choose_req_valids[6] <= (soc_videosoc_sdram_bankmachine6_cmd_valid & ((soc_videosoc_sdram_bankmachine6_cmd_payload_is_cmd & soc_videosoc_sdram_choose_req_want_cmds) | ((soc_videosoc_sdram_bankmachine6_cmd_payload_is_read == soc_videosoc_sdram_choose_req_want_reads) & (soc_videosoc_sdram_bankmachine6_cmd_payload_is_write == soc_videosoc_sdram_choose_req_want_writes))));
	soc_videosoc_sdram_choose_req_valids[7] <= (soc_videosoc_sdram_bankmachine7_cmd_valid & ((soc_videosoc_sdram_bankmachine7_cmd_payload_is_cmd & soc_videosoc_sdram_choose_req_want_cmds) | ((soc_videosoc_sdram_bankmachine7_cmd_payload_is_read == soc_videosoc_sdram_choose_req_want_reads) & (soc_videosoc_sdram_bankmachine7_cmd_payload_is_write == soc_videosoc_sdram_choose_req_want_writes))));
end
assign soc_videosoc_sdram_choose_req_request = soc_videosoc_sdram_choose_req_valids;
assign soc_videosoc_sdram_choose_req_cmd_valid = vns_comb_rhs_array_muxed6;
assign soc_videosoc_sdram_choose_req_cmd_payload_a = vns_comb_rhs_array_muxed7;
assign soc_videosoc_sdram_choose_req_cmd_payload_ba = vns_comb_rhs_array_muxed8;
assign soc_videosoc_sdram_choose_req_cmd_payload_is_read = vns_comb_rhs_array_muxed9;
assign soc_videosoc_sdram_choose_req_cmd_payload_is_write = vns_comb_rhs_array_muxed10;
assign soc_videosoc_sdram_choose_req_cmd_payload_is_cmd = vns_comb_rhs_array_muxed11;
always @(*) begin
	soc_videosoc_sdram_choose_req_cmd_payload_cas <= 1'd0;
	if (soc_videosoc_sdram_choose_req_cmd_valid) begin
		soc_videosoc_sdram_choose_req_cmd_payload_cas <= vns_comb_t_array_muxed3;
	end
end
always @(*) begin
	soc_videosoc_sdram_choose_req_cmd_payload_ras <= 1'd0;
	if (soc_videosoc_sdram_choose_req_cmd_valid) begin
		soc_videosoc_sdram_choose_req_cmd_payload_ras <= vns_comb_t_array_muxed4;
	end
end
always @(*) begin
	soc_videosoc_sdram_choose_req_cmd_payload_we <= 1'd0;
	if (soc_videosoc_sdram_choose_req_cmd_valid) begin
		soc_videosoc_sdram_choose_req_cmd_payload_we <= vns_comb_t_array_muxed5;
	end
end
always @(*) begin
	soc_videosoc_sdram_bankmachine0_cmd_ready <= 1'd0;
	if (((soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_ready) & (soc_videosoc_sdram_choose_cmd_grant == 1'd0))) begin
		soc_videosoc_sdram_bankmachine0_cmd_ready <= 1'd1;
	end
	if (((soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_ready) & (soc_videosoc_sdram_choose_req_grant == 1'd0))) begin
		soc_videosoc_sdram_bankmachine0_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	soc_videosoc_sdram_bankmachine1_cmd_ready <= 1'd0;
	if (((soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_ready) & (soc_videosoc_sdram_choose_cmd_grant == 1'd1))) begin
		soc_videosoc_sdram_bankmachine1_cmd_ready <= 1'd1;
	end
	if (((soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_ready) & (soc_videosoc_sdram_choose_req_grant == 1'd1))) begin
		soc_videosoc_sdram_bankmachine1_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	soc_videosoc_sdram_bankmachine2_cmd_ready <= 1'd0;
	if (((soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_ready) & (soc_videosoc_sdram_choose_cmd_grant == 2'd2))) begin
		soc_videosoc_sdram_bankmachine2_cmd_ready <= 1'd1;
	end
	if (((soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_ready) & (soc_videosoc_sdram_choose_req_grant == 2'd2))) begin
		soc_videosoc_sdram_bankmachine2_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	soc_videosoc_sdram_bankmachine3_cmd_ready <= 1'd0;
	if (((soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_ready) & (soc_videosoc_sdram_choose_cmd_grant == 2'd3))) begin
		soc_videosoc_sdram_bankmachine3_cmd_ready <= 1'd1;
	end
	if (((soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_ready) & (soc_videosoc_sdram_choose_req_grant == 2'd3))) begin
		soc_videosoc_sdram_bankmachine3_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	soc_videosoc_sdram_bankmachine4_cmd_ready <= 1'd0;
	if (((soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_ready) & (soc_videosoc_sdram_choose_cmd_grant == 3'd4))) begin
		soc_videosoc_sdram_bankmachine4_cmd_ready <= 1'd1;
	end
	if (((soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_ready) & (soc_videosoc_sdram_choose_req_grant == 3'd4))) begin
		soc_videosoc_sdram_bankmachine4_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	soc_videosoc_sdram_bankmachine5_cmd_ready <= 1'd0;
	if (((soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_ready) & (soc_videosoc_sdram_choose_cmd_grant == 3'd5))) begin
		soc_videosoc_sdram_bankmachine5_cmd_ready <= 1'd1;
	end
	if (((soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_ready) & (soc_videosoc_sdram_choose_req_grant == 3'd5))) begin
		soc_videosoc_sdram_bankmachine5_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	soc_videosoc_sdram_bankmachine6_cmd_ready <= 1'd0;
	if (((soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_ready) & (soc_videosoc_sdram_choose_cmd_grant == 3'd6))) begin
		soc_videosoc_sdram_bankmachine6_cmd_ready <= 1'd1;
	end
	if (((soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_ready) & (soc_videosoc_sdram_choose_req_grant == 3'd6))) begin
		soc_videosoc_sdram_bankmachine6_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	soc_videosoc_sdram_bankmachine7_cmd_ready <= 1'd0;
	if (((soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_ready) & (soc_videosoc_sdram_choose_cmd_grant == 3'd7))) begin
		soc_videosoc_sdram_bankmachine7_cmd_ready <= 1'd1;
	end
	if (((soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_ready) & (soc_videosoc_sdram_choose_req_grant == 3'd7))) begin
		soc_videosoc_sdram_bankmachine7_cmd_ready <= 1'd1;
	end
end
assign soc_videosoc_sdram_choose_req_ce = soc_videosoc_sdram_choose_req_cmd_ready;
assign soc_videosoc_sdram_dfi_p0_cke = 1'd1;
assign soc_videosoc_sdram_dfi_p0_cs_n = 1'd0;
assign soc_videosoc_sdram_dfi_p0_odt = 1'd1;
assign soc_videosoc_sdram_dfi_p0_reset_n = 1'd1;
assign soc_videosoc_sdram_dfi_p1_cke = 1'd1;
assign soc_videosoc_sdram_dfi_p1_cs_n = 1'd0;
assign soc_videosoc_sdram_dfi_p1_odt = 1'd1;
assign soc_videosoc_sdram_dfi_p1_reset_n = 1'd1;
assign soc_videosoc_sdram_dfi_p2_cke = 1'd1;
assign soc_videosoc_sdram_dfi_p2_cs_n = 1'd0;
assign soc_videosoc_sdram_dfi_p2_odt = 1'd1;
assign soc_videosoc_sdram_dfi_p2_reset_n = 1'd1;
assign soc_videosoc_sdram_dfi_p3_cke = 1'd1;
assign soc_videosoc_sdram_dfi_p3_cs_n = 1'd0;
assign soc_videosoc_sdram_dfi_p3_odt = 1'd1;
assign soc_videosoc_sdram_dfi_p3_reset_n = 1'd1;
always @(*) begin
	soc_videosoc_sdram_en1 <= 1'd0;
	soc_videosoc_sdram_choose_req_cmd_ready <= 1'd0;
	soc_videosoc_sdram_cmd_ready <= 1'd0;
	vns_multiplexer_next_state <= 4'd0;
	soc_videosoc_sdram_sel0 <= 2'd0;
	soc_videosoc_sdram_choose_cmd_cmd_ready <= 1'd0;
	soc_videosoc_sdram_sel1 <= 2'd0;
	soc_videosoc_sdram_en0 <= 1'd0;
	soc_videosoc_sdram_sel2 <= 2'd0;
	soc_videosoc_sdram_sel3 <= 2'd0;
	soc_videosoc_sdram_choose_req_want_reads <= 1'd0;
	soc_videosoc_sdram_choose_req_want_writes <= 1'd0;
	vns_multiplexer_next_state <= vns_multiplexer_state;
	case (vns_multiplexer_state)
		1'd1: begin
			soc_videosoc_sdram_en1 <= 1'd1;
			soc_videosoc_sdram_choose_req_want_writes <= 1'd1;
			soc_videosoc_sdram_choose_cmd_cmd_ready <= 1'd1;
			soc_videosoc_sdram_choose_req_cmd_ready <= 1'd1;
			soc_videosoc_sdram_sel0 <= 1'd1;
			soc_videosoc_sdram_sel1 <= 1'd0;
			soc_videosoc_sdram_sel2 <= 2'd2;
			soc_videosoc_sdram_sel3 <= 1'd0;
			if (soc_videosoc_sdram_read_available) begin
				if (((~soc_videosoc_sdram_write_available) | soc_videosoc_sdram_max_time1)) begin
					vns_multiplexer_next_state <= 4'd8;
				end
			end
			if (soc_videosoc_sdram_go_to_refresh) begin
				vns_multiplexer_next_state <= 2'd2;
			end
		end
		2'd2: begin
			soc_videosoc_sdram_sel0 <= 2'd3;
			soc_videosoc_sdram_cmd_ready <= 1'd1;
			if (soc_videosoc_sdram_cmd_last) begin
				vns_multiplexer_next_state <= 1'd0;
			end
		end
		2'd3: begin
			vns_multiplexer_next_state <= 3'd4;
		end
		3'd4: begin
			vns_multiplexer_next_state <= 3'd5;
		end
		3'd5: begin
			vns_multiplexer_next_state <= 3'd6;
		end
		3'd6: begin
			vns_multiplexer_next_state <= 3'd7;
		end
		3'd7: begin
			vns_multiplexer_next_state <= 1'd1;
		end
		4'd8: begin
			vns_multiplexer_next_state <= 4'd9;
		end
		4'd9: begin
			vns_multiplexer_next_state <= 4'd10;
		end
		4'd10: begin
			vns_multiplexer_next_state <= 4'd11;
		end
		4'd11: begin
			vns_multiplexer_next_state <= 4'd12;
		end
		4'd12: begin
			vns_multiplexer_next_state <= 4'd13;
		end
		4'd13: begin
			vns_multiplexer_next_state <= 4'd14;
		end
		4'd14: begin
			vns_multiplexer_next_state <= 1'd0;
		end
		default: begin
			soc_videosoc_sdram_en0 <= 1'd1;
			soc_videosoc_sdram_choose_req_want_reads <= 1'd1;
			soc_videosoc_sdram_choose_cmd_cmd_ready <= 1'd1;
			soc_videosoc_sdram_choose_req_cmd_ready <= 1'd1;
			soc_videosoc_sdram_sel0 <= 2'd2;
			soc_videosoc_sdram_sel1 <= 1'd1;
			soc_videosoc_sdram_sel2 <= 1'd0;
			soc_videosoc_sdram_sel3 <= 1'd0;
			if (soc_videosoc_sdram_write_available) begin
				if (((~soc_videosoc_sdram_read_available) | soc_videosoc_sdram_max_time0)) begin
					vns_multiplexer_next_state <= 2'd3;
				end
			end
			if (soc_videosoc_sdram_go_to_refresh) begin
				vns_multiplexer_next_state <= 2'd2;
			end
		end
	endcase
end
assign vns_cba0 = soc_videosoc_port_cmd_payload_adr[9:7];
assign vns_rca0 = {soc_videosoc_port_cmd_payload_adr[24:10], soc_videosoc_port_cmd_payload_adr[6:0]};
assign vns_cba1 = soc_litedramcrossbar_cmd_payload_adr[9:7];
assign vns_rca1 = {soc_litedramcrossbar_cmd_payload_adr[24:10], soc_litedramcrossbar_cmd_payload_adr[6:0]};
assign vns_cba2 = soc_hdmi_out0_dram_port_cmd_payload_adr[9:7];
assign vns_rca2 = {soc_hdmi_out0_dram_port_cmd_payload_adr[24:10], soc_hdmi_out0_dram_port_cmd_payload_adr[6:0]};
assign vns_roundrobin0_request = {(((vns_cba2 == 1'd0) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid), (((vns_cba1 == 1'd0) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid), (((vns_cba0 == 1'd0) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videosoc_port_cmd_valid)};
assign vns_roundrobin0_ce = ((~soc_videosoc_sdram_interface_bank0_valid) & (~soc_videosoc_sdram_interface_bank0_lock));
assign soc_videosoc_sdram_interface_bank0_adr = vns_comb_rhs_array_muxed12;
assign soc_videosoc_sdram_interface_bank0_we = vns_comb_rhs_array_muxed13;
assign soc_videosoc_sdram_interface_bank0_valid = vns_comb_rhs_array_muxed14;
assign vns_roundrobin1_request = {(((vns_cba2 == 1'd1) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid), (((vns_cba1 == 1'd1) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid), (((vns_cba0 == 1'd1) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videosoc_port_cmd_valid)};
assign vns_roundrobin1_ce = ((~soc_videosoc_sdram_interface_bank1_valid) & (~soc_videosoc_sdram_interface_bank1_lock));
assign soc_videosoc_sdram_interface_bank1_adr = vns_comb_rhs_array_muxed15;
assign soc_videosoc_sdram_interface_bank1_we = vns_comb_rhs_array_muxed16;
assign soc_videosoc_sdram_interface_bank1_valid = vns_comb_rhs_array_muxed17;
assign vns_roundrobin2_request = {(((vns_cba2 == 2'd2) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid), (((vns_cba1 == 2'd2) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid), (((vns_cba0 == 2'd2) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videosoc_port_cmd_valid)};
assign vns_roundrobin2_ce = ((~soc_videosoc_sdram_interface_bank2_valid) & (~soc_videosoc_sdram_interface_bank2_lock));
assign soc_videosoc_sdram_interface_bank2_adr = vns_comb_rhs_array_muxed18;
assign soc_videosoc_sdram_interface_bank2_we = vns_comb_rhs_array_muxed19;
assign soc_videosoc_sdram_interface_bank2_valid = vns_comb_rhs_array_muxed20;
assign vns_roundrobin3_request = {(((vns_cba2 == 2'd3) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid), (((vns_cba1 == 2'd3) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid), (((vns_cba0 == 2'd3) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videosoc_port_cmd_valid)};
assign vns_roundrobin3_ce = ((~soc_videosoc_sdram_interface_bank3_valid) & (~soc_videosoc_sdram_interface_bank3_lock));
assign soc_videosoc_sdram_interface_bank3_adr = vns_comb_rhs_array_muxed21;
assign soc_videosoc_sdram_interface_bank3_we = vns_comb_rhs_array_muxed22;
assign soc_videosoc_sdram_interface_bank3_valid = vns_comb_rhs_array_muxed23;
assign vns_roundrobin4_request = {(((vns_cba2 == 3'd4) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid), (((vns_cba1 == 3'd4) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid), (((vns_cba0 == 3'd4) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videosoc_port_cmd_valid)};
assign vns_roundrobin4_ce = ((~soc_videosoc_sdram_interface_bank4_valid) & (~soc_videosoc_sdram_interface_bank4_lock));
assign soc_videosoc_sdram_interface_bank4_adr = vns_comb_rhs_array_muxed24;
assign soc_videosoc_sdram_interface_bank4_we = vns_comb_rhs_array_muxed25;
assign soc_videosoc_sdram_interface_bank4_valid = vns_comb_rhs_array_muxed26;
assign vns_roundrobin5_request = {(((vns_cba2 == 3'd5) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid), (((vns_cba1 == 3'd5) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid), (((vns_cba0 == 3'd5) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videosoc_port_cmd_valid)};
assign vns_roundrobin5_ce = ((~soc_videosoc_sdram_interface_bank5_valid) & (~soc_videosoc_sdram_interface_bank5_lock));
assign soc_videosoc_sdram_interface_bank5_adr = vns_comb_rhs_array_muxed27;
assign soc_videosoc_sdram_interface_bank5_we = vns_comb_rhs_array_muxed28;
assign soc_videosoc_sdram_interface_bank5_valid = vns_comb_rhs_array_muxed29;
assign vns_roundrobin6_request = {(((vns_cba2 == 3'd6) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid), (((vns_cba1 == 3'd6) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid), (((vns_cba0 == 3'd6) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videosoc_port_cmd_valid)};
assign vns_roundrobin6_ce = ((~soc_videosoc_sdram_interface_bank6_valid) & (~soc_videosoc_sdram_interface_bank6_lock));
assign soc_videosoc_sdram_interface_bank6_adr = vns_comb_rhs_array_muxed30;
assign soc_videosoc_sdram_interface_bank6_we = vns_comb_rhs_array_muxed31;
assign soc_videosoc_sdram_interface_bank6_valid = vns_comb_rhs_array_muxed32;
assign vns_roundrobin7_request = {(((vns_cba2 == 3'd7) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid), (((vns_cba1 == 3'd7) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid), (((vns_cba0 == 3'd7) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))))) & soc_videosoc_port_cmd_valid)};
assign vns_roundrobin7_ce = ((~soc_videosoc_sdram_interface_bank7_valid) & (~soc_videosoc_sdram_interface_bank7_lock));
assign soc_videosoc_sdram_interface_bank7_adr = vns_comb_rhs_array_muxed33;
assign soc_videosoc_sdram_interface_bank7_we = vns_comb_rhs_array_muxed34;
assign soc_videosoc_sdram_interface_bank7_valid = vns_comb_rhs_array_muxed35;
assign soc_videosoc_port_cmd_ready = ((((((((1'd0 | (((vns_roundrobin0_grant == 1'd0) & ((vns_cba0 == 1'd0) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0)))))) & soc_videosoc_sdram_interface_bank0_ready)) | (((vns_roundrobin1_grant == 1'd0) & ((vns_cba0 == 1'd1) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0)))))) & soc_videosoc_sdram_interface_bank1_ready)) | (((vns_roundrobin2_grant == 1'd0) & ((vns_cba0 == 2'd2) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0)))))) & soc_videosoc_sdram_interface_bank2_ready)) | (((vns_roundrobin3_grant == 1'd0) & ((vns_cba0 == 2'd3) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0)))))) & soc_videosoc_sdram_interface_bank3_ready)) | (((vns_roundrobin4_grant == 1'd0) & ((vns_cba0 == 3'd4) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0)))))) & soc_videosoc_sdram_interface_bank4_ready)) | (((vns_roundrobin5_grant == 1'd0) & ((vns_cba0 == 3'd5) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0)))))) & soc_videosoc_sdram_interface_bank5_ready)) | (((vns_roundrobin6_grant == 1'd0) & ((vns_cba0 == 3'd6) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0)))))) & soc_videosoc_sdram_interface_bank6_ready)) | (((vns_roundrobin7_grant == 1'd0) & ((vns_cba0 == 3'd7) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0)))))) & soc_videosoc_sdram_interface_bank7_ready));
assign soc_litedramcrossbar_cmd_ready = ((((((((1'd0 | (((vns_roundrobin0_grant == 1'd1) & ((vns_cba1 == 1'd0) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1)))))) & soc_videosoc_sdram_interface_bank0_ready)) | (((vns_roundrobin1_grant == 1'd1) & ((vns_cba1 == 1'd1) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1)))))) & soc_videosoc_sdram_interface_bank1_ready)) | (((vns_roundrobin2_grant == 1'd1) & ((vns_cba1 == 2'd2) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1)))))) & soc_videosoc_sdram_interface_bank2_ready)) | (((vns_roundrobin3_grant == 1'd1) & ((vns_cba1 == 2'd3) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1)))))) & soc_videosoc_sdram_interface_bank3_ready)) | (((vns_roundrobin4_grant == 1'd1) & ((vns_cba1 == 3'd4) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1)))))) & soc_videosoc_sdram_interface_bank4_ready)) | (((vns_roundrobin5_grant == 1'd1) & ((vns_cba1 == 3'd5) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1)))))) & soc_videosoc_sdram_interface_bank5_ready)) | (((vns_roundrobin6_grant == 1'd1) & ((vns_cba1 == 3'd6) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1)))))) & soc_videosoc_sdram_interface_bank6_ready)) | (((vns_roundrobin7_grant == 1'd1) & ((vns_cba1 == 3'd7) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1)))))) & soc_videosoc_sdram_interface_bank7_ready));
assign soc_hdmi_out0_dram_port_cmd_ready = ((((((((1'd0 | (((vns_roundrobin0_grant == 2'd2) & ((vns_cba2 == 1'd0) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2)))))) & soc_videosoc_sdram_interface_bank0_ready)) | (((vns_roundrobin1_grant == 2'd2) & ((vns_cba2 == 1'd1) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2)))))) & soc_videosoc_sdram_interface_bank1_ready)) | (((vns_roundrobin2_grant == 2'd2) & ((vns_cba2 == 2'd2) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2)))))) & soc_videosoc_sdram_interface_bank2_ready)) | (((vns_roundrobin3_grant == 2'd2) & ((vns_cba2 == 2'd3) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2)))))) & soc_videosoc_sdram_interface_bank3_ready)) | (((vns_roundrobin4_grant == 2'd2) & ((vns_cba2 == 3'd4) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2)))))) & soc_videosoc_sdram_interface_bank4_ready)) | (((vns_roundrobin5_grant == 2'd2) & ((vns_cba2 == 3'd5) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2)))))) & soc_videosoc_sdram_interface_bank5_ready)) | (((vns_roundrobin6_grant == 2'd2) & ((vns_cba2 == 3'd6) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2)))))) & soc_videosoc_sdram_interface_bank6_ready)) | (((vns_roundrobin7_grant == 2'd2) & ((vns_cba2 == 3'd7) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2)))))) & soc_videosoc_sdram_interface_bank7_ready));
assign soc_videosoc_port_wdata_ready = vns_new_master_wdata_ready2;
assign soc_litedramcrossbar_wdata_ready = vns_new_master_wdata_ready5;
assign soc_hdmi_out0_dram_port_wdata_ready = vns_new_master_wdata_ready8;
assign soc_videosoc_port_rdata_valid = vns_new_master_rdata_valid6;
assign soc_litedramcrossbar_rdata_valid = vns_new_master_rdata_valid13;
assign soc_hdmi_out0_dram_port_rdata_valid = vns_new_master_rdata_valid20;
always @(*) begin
	soc_videosoc_sdram_interface_wdata_we <= 16'd0;
	soc_videosoc_sdram_interface_wdata <= 128'd0;
	case ({vns_new_master_wdata_ready8, vns_new_master_wdata_ready5, vns_new_master_wdata_ready2})
		1'd1: begin
			soc_videosoc_sdram_interface_wdata <= soc_videosoc_port_wdata_payload_data;
			soc_videosoc_sdram_interface_wdata_we <= soc_videosoc_port_wdata_payload_we;
		end
		2'd2: begin
			soc_videosoc_sdram_interface_wdata <= soc_litedramcrossbar_wdata_payload_data;
			soc_videosoc_sdram_interface_wdata_we <= soc_litedramcrossbar_wdata_payload_we;
		end
		3'd4: begin
			soc_videosoc_sdram_interface_wdata <= soc_hdmi_out0_dram_port_wdata_payload_data;
			soc_videosoc_sdram_interface_wdata_we <= soc_hdmi_out0_dram_port_wdata_payload_we;
		end
		default: begin
			soc_videosoc_sdram_interface_wdata <= 1'd0;
			soc_videosoc_sdram_interface_wdata_we <= 1'd0;
		end
	endcase
end
assign soc_videosoc_port_rdata_payload_data = soc_videosoc_sdram_interface_rdata;
assign soc_litedramcrossbar_rdata_payload_data = soc_videosoc_sdram_interface_rdata;
assign soc_hdmi_out0_dram_port_rdata_payload_data = soc_videosoc_sdram_interface_rdata;
assign soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_din = {soc_hdmi_out0_dram_port_cmd_fifo_fifo_in_last, soc_hdmi_out0_dram_port_cmd_fifo_fifo_in_first, soc_hdmi_out0_dram_port_cmd_fifo_fifo_in_payload_adr, soc_hdmi_out0_dram_port_cmd_fifo_fifo_in_payload_we};
assign {soc_hdmi_out0_dram_port_cmd_fifo_fifo_out_last, soc_hdmi_out0_dram_port_cmd_fifo_fifo_out_first, soc_hdmi_out0_dram_port_cmd_fifo_fifo_out_payload_adr, soc_hdmi_out0_dram_port_cmd_fifo_fifo_out_payload_we} = soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_dout;
assign soc_hdmi_out0_dram_port_cmd_fifo_sink_ready = soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_writable;
assign soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_we = soc_hdmi_out0_dram_port_cmd_fifo_sink_valid;
assign soc_hdmi_out0_dram_port_cmd_fifo_fifo_in_first = soc_hdmi_out0_dram_port_cmd_fifo_sink_first;
assign soc_hdmi_out0_dram_port_cmd_fifo_fifo_in_last = soc_hdmi_out0_dram_port_cmd_fifo_sink_last;
assign soc_hdmi_out0_dram_port_cmd_fifo_fifo_in_payload_we = soc_hdmi_out0_dram_port_cmd_fifo_sink_payload_we;
assign soc_hdmi_out0_dram_port_cmd_fifo_fifo_in_payload_adr = soc_hdmi_out0_dram_port_cmd_fifo_sink_payload_adr;
assign soc_hdmi_out0_dram_port_cmd_fifo_source_valid = soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_readable;
assign soc_hdmi_out0_dram_port_cmd_fifo_source_first = soc_hdmi_out0_dram_port_cmd_fifo_fifo_out_first;
assign soc_hdmi_out0_dram_port_cmd_fifo_source_last = soc_hdmi_out0_dram_port_cmd_fifo_fifo_out_last;
assign soc_hdmi_out0_dram_port_cmd_fifo_source_payload_we = soc_hdmi_out0_dram_port_cmd_fifo_fifo_out_payload_we;
assign soc_hdmi_out0_dram_port_cmd_fifo_source_payload_adr = soc_hdmi_out0_dram_port_cmd_fifo_fifo_out_payload_adr;
assign soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_re = soc_hdmi_out0_dram_port_cmd_fifo_source_ready;
assign soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_ce = (soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_writable & soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_we);
assign soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_ce = (soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_readable & soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_re);
assign soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_writable = (((soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q[2] == soc_hdmi_out0_dram_port_cmd_fifo_consume_wdomain[2]) | (soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q[1] == soc_hdmi_out0_dram_port_cmd_fifo_consume_wdomain[1])) | (soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q[0] != soc_hdmi_out0_dram_port_cmd_fifo_consume_wdomain[0]));
assign soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_readable = (soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q != soc_hdmi_out0_dram_port_cmd_fifo_produce_rdomain);
assign soc_hdmi_out0_dram_port_cmd_fifo_wrport_adr = soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_binary[1:0];
assign soc_hdmi_out0_dram_port_cmd_fifo_wrport_dat_w = soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_din;
assign soc_hdmi_out0_dram_port_cmd_fifo_wrport_we = soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_ce;
assign soc_hdmi_out0_dram_port_cmd_fifo_rdport_adr = soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary[1:0];
assign soc_hdmi_out0_dram_port_cmd_fifo_asyncfifo_dout = soc_hdmi_out0_dram_port_cmd_fifo_rdport_dat_r;
always @(*) begin
	soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next_binary <= 3'd0;
	if (soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_ce) begin
		soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next_binary <= (soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_binary + 1'd1);
	end else begin
		soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next_binary <= soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_binary;
	end
end
assign soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next = (soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next_binary ^ soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next_binary[2:1]);
always @(*) begin
	soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary <= 3'd0;
	if (soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_ce) begin
		soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary <= (soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_binary + 1'd1);
	end else begin
		soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary <= soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_binary;
	end
end
assign soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next = (soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary ^ soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary[2:1]);
assign soc_hdmi_out0_dram_port_cmd_fifo_sink_valid = soc_hdmi_out0_dram_port_litedramport0_cmd_valid;
assign soc_hdmi_out0_dram_port_litedramport0_cmd_ready = soc_hdmi_out0_dram_port_cmd_fifo_sink_ready;
assign soc_hdmi_out0_dram_port_cmd_fifo_sink_first = soc_hdmi_out0_dram_port_litedramport0_cmd_first;
assign soc_hdmi_out0_dram_port_cmd_fifo_sink_last = soc_hdmi_out0_dram_port_litedramport0_cmd_last;
assign soc_hdmi_out0_dram_port_cmd_fifo_sink_payload_we = soc_hdmi_out0_dram_port_litedramport0_cmd_payload_we;
assign soc_hdmi_out0_dram_port_cmd_fifo_sink_payload_adr = soc_hdmi_out0_dram_port_litedramport0_cmd_payload_adr;
assign soc_hdmi_out0_dram_port_cmd_valid = soc_hdmi_out0_dram_port_cmd_fifo_source_valid;
assign soc_hdmi_out0_dram_port_cmd_fifo_source_ready = soc_hdmi_out0_dram_port_cmd_ready;
assign soc_hdmi_out0_dram_port_cmd_first = soc_hdmi_out0_dram_port_cmd_fifo_source_first;
assign soc_hdmi_out0_dram_port_cmd_last = soc_hdmi_out0_dram_port_cmd_fifo_source_last;
assign soc_hdmi_out0_dram_port_cmd_payload_we = soc_hdmi_out0_dram_port_cmd_fifo_source_payload_we;
assign soc_hdmi_out0_dram_port_cmd_payload_adr = soc_hdmi_out0_dram_port_cmd_fifo_source_payload_adr;
assign soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_din = {soc_hdmi_out0_dram_port_rdata_fifo_fifo_in_last, soc_hdmi_out0_dram_port_rdata_fifo_fifo_in_first, soc_hdmi_out0_dram_port_rdata_fifo_fifo_in_payload_data};
assign {soc_hdmi_out0_dram_port_rdata_fifo_fifo_out_last, soc_hdmi_out0_dram_port_rdata_fifo_fifo_out_first, soc_hdmi_out0_dram_port_rdata_fifo_fifo_out_payload_data} = soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_dout;
assign soc_hdmi_out0_dram_port_rdata_fifo_sink_ready = soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_writable;
assign soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_we = soc_hdmi_out0_dram_port_rdata_fifo_sink_valid;
assign soc_hdmi_out0_dram_port_rdata_fifo_fifo_in_first = soc_hdmi_out0_dram_port_rdata_fifo_sink_first;
assign soc_hdmi_out0_dram_port_rdata_fifo_fifo_in_last = soc_hdmi_out0_dram_port_rdata_fifo_sink_last;
assign soc_hdmi_out0_dram_port_rdata_fifo_fifo_in_payload_data = soc_hdmi_out0_dram_port_rdata_fifo_sink_payload_data;
assign soc_hdmi_out0_dram_port_rdata_fifo_source_valid = soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_readable;
assign soc_hdmi_out0_dram_port_rdata_fifo_source_first = soc_hdmi_out0_dram_port_rdata_fifo_fifo_out_first;
assign soc_hdmi_out0_dram_port_rdata_fifo_source_last = soc_hdmi_out0_dram_port_rdata_fifo_fifo_out_last;
assign soc_hdmi_out0_dram_port_rdata_fifo_source_payload_data = soc_hdmi_out0_dram_port_rdata_fifo_fifo_out_payload_data;
assign soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_re = soc_hdmi_out0_dram_port_rdata_fifo_source_ready;
assign soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_ce = (soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_writable & soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_we);
assign soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_ce = (soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_readable & soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_re);
assign soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_writable = (((soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q[4] == soc_hdmi_out0_dram_port_rdata_fifo_consume_wdomain[4]) | (soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q[3] == soc_hdmi_out0_dram_port_rdata_fifo_consume_wdomain[3])) | (soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q[2:0] != soc_hdmi_out0_dram_port_rdata_fifo_consume_wdomain[2:0]));
assign soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_readable = (soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q != soc_hdmi_out0_dram_port_rdata_fifo_produce_rdomain);
assign soc_hdmi_out0_dram_port_rdata_fifo_wrport_adr = soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_binary[3:0];
assign soc_hdmi_out0_dram_port_rdata_fifo_wrport_dat_w = soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_din;
assign soc_hdmi_out0_dram_port_rdata_fifo_wrport_we = soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_ce;
assign soc_hdmi_out0_dram_port_rdata_fifo_rdport_adr = soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary[3:0];
assign soc_hdmi_out0_dram_port_rdata_fifo_asyncfifo_dout = soc_hdmi_out0_dram_port_rdata_fifo_rdport_dat_r;
always @(*) begin
	soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next_binary <= 5'd0;
	if (soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_ce) begin
		soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next_binary <= (soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_binary + 1'd1);
	end else begin
		soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next_binary <= soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_binary;
	end
end
assign soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next = (soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next_binary ^ soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next_binary[4:1]);
always @(*) begin
	soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary <= 5'd0;
	if (soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_ce) begin
		soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary <= (soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_binary + 1'd1);
	end else begin
		soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary <= soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_binary;
	end
end
assign soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next = (soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary ^ soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary[4:1]);
assign soc_hdmi_out0_dram_port_rdata_fifo_sink_valid = soc_hdmi_out0_dram_port_rdata_valid;
assign soc_hdmi_out0_dram_port_rdata_ready = soc_hdmi_out0_dram_port_rdata_fifo_sink_ready;
assign soc_hdmi_out0_dram_port_rdata_fifo_sink_first = soc_hdmi_out0_dram_port_rdata_first;
assign soc_hdmi_out0_dram_port_rdata_fifo_sink_last = soc_hdmi_out0_dram_port_rdata_last;
assign soc_hdmi_out0_dram_port_rdata_fifo_sink_payload_data = soc_hdmi_out0_dram_port_rdata_payload_data;
assign soc_hdmi_out0_dram_port_litedramport0_rdata_valid = soc_hdmi_out0_dram_port_rdata_fifo_source_valid;
assign soc_hdmi_out0_dram_port_rdata_fifo_source_ready = soc_hdmi_out0_dram_port_litedramport0_rdata_ready;
assign soc_hdmi_out0_dram_port_litedramport0_rdata_first = soc_hdmi_out0_dram_port_rdata_fifo_source_first;
assign soc_hdmi_out0_dram_port_litedramport0_rdata_last = soc_hdmi_out0_dram_port_rdata_fifo_source_last;
assign soc_hdmi_out0_dram_port_litedramport0_rdata_payload_data = soc_hdmi_out0_dram_port_rdata_fifo_source_payload_data;
always @(*) begin
	soc_hdmi_out0_dram_port_litedramport0_cmd_valid <= 1'd0;
	soc_hdmi_out0_dram_port_litedramport1_cmd_ready <= 1'd0;
	soc_hdmi_out0_dram_port_litedramport0_cmd_payload_adr <= 25'd0;
	soc_hdmi_out0_dram_port_counter_ce <= 1'd0;
	if (soc_hdmi_out0_dram_port_litedramport1_cmd_valid) begin
		if ((soc_hdmi_out0_dram_port_counter == 1'd0)) begin
			soc_hdmi_out0_dram_port_litedramport0_cmd_valid <= 1'd1;
			soc_hdmi_out0_dram_port_litedramport0_cmd_payload_adr <= soc_hdmi_out0_dram_port_litedramport1_cmd_payload_adr[27:3];
			soc_hdmi_out0_dram_port_litedramport1_cmd_ready <= soc_hdmi_out0_dram_port_litedramport0_cmd_ready;
			soc_hdmi_out0_dram_port_counter_ce <= soc_hdmi_out0_dram_port_litedramport0_cmd_ready;
		end else begin
			soc_hdmi_out0_dram_port_litedramport1_cmd_ready <= 1'd1;
			soc_hdmi_out0_dram_port_counter_ce <= 1'd1;
		end
	end
end
always @(*) begin
	soc_hdmi_out0_dram_port_cmd_buffer_sink_valid <= 1'd0;
	soc_hdmi_out0_dram_port_cmd_buffer_sink_payload_sel <= 8'd0;
	if ((soc_hdmi_out0_dram_port_litedramport0_cmd_valid & soc_hdmi_out0_dram_port_litedramport0_cmd_ready)) begin
		soc_hdmi_out0_dram_port_cmd_buffer_sink_valid <= 1'd1;
		soc_hdmi_out0_dram_port_cmd_buffer_sink_payload_sel <= 8'd255;
	end
end
assign soc_hdmi_out0_dram_port_rdata_buffer_sink_valid = soc_hdmi_out0_dram_port_litedramport0_rdata_valid;
assign soc_hdmi_out0_dram_port_litedramport0_rdata_ready = soc_hdmi_out0_dram_port_rdata_buffer_sink_ready;
assign soc_hdmi_out0_dram_port_rdata_buffer_sink_first = soc_hdmi_out0_dram_port_litedramport0_rdata_first;
assign soc_hdmi_out0_dram_port_rdata_buffer_sink_last = soc_hdmi_out0_dram_port_litedramport0_rdata_last;
assign soc_hdmi_out0_dram_port_rdata_buffer_sink_payload_data = soc_hdmi_out0_dram_port_litedramport0_rdata_payload_data;
assign soc_hdmi_out0_dram_port_rdata_converter_sink_valid = soc_hdmi_out0_dram_port_rdata_buffer_source_valid;
assign soc_hdmi_out0_dram_port_rdata_buffer_source_ready = soc_hdmi_out0_dram_port_rdata_converter_sink_ready;
assign soc_hdmi_out0_dram_port_rdata_converter_sink_first = soc_hdmi_out0_dram_port_rdata_buffer_source_first;
assign soc_hdmi_out0_dram_port_rdata_converter_sink_last = soc_hdmi_out0_dram_port_rdata_buffer_source_last;
assign soc_hdmi_out0_dram_port_rdata_converter_sink_payload_data = soc_hdmi_out0_dram_port_rdata_buffer_source_payload_data;
assign soc_hdmi_out0_dram_port_rdata_chunk_valid = ((soc_hdmi_out0_dram_port_cmd_buffer_source_payload_sel & soc_hdmi_out0_dram_port_rdata_chunk) != 1'd0);
always @(*) begin
	soc_hdmi_out0_dram_port_litedramport1_rdata_valid <= 1'd0;
	soc_hdmi_out0_dram_port_rdata_converter_source_ready <= 1'd0;
	soc_hdmi_out0_dram_port_litedramport1_rdata_payload_data <= 16'd0;
	if (soc_hdmi_out0_dram_port_litedramport1_flush) begin
		soc_hdmi_out0_dram_port_rdata_converter_source_ready <= 1'd1;
	end else begin
		if (soc_hdmi_out0_dram_port_cmd_buffer_source_valid) begin
			if (soc_hdmi_out0_dram_port_rdata_chunk_valid) begin
				soc_hdmi_out0_dram_port_litedramport1_rdata_valid <= soc_hdmi_out0_dram_port_rdata_converter_source_valid;
				soc_hdmi_out0_dram_port_litedramport1_rdata_payload_data <= soc_hdmi_out0_dram_port_rdata_converter_source_payload_data;
				soc_hdmi_out0_dram_port_rdata_converter_source_ready <= soc_hdmi_out0_dram_port_litedramport1_rdata_ready;
			end else begin
				soc_hdmi_out0_dram_port_rdata_converter_source_ready <= 1'd1;
			end
		end
	end
end
assign soc_hdmi_out0_dram_port_cmd_buffer_source_ready = (soc_hdmi_out0_dram_port_rdata_converter_source_ready & soc_hdmi_out0_dram_port_rdata_chunk[7]);
assign soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_din = {soc_hdmi_out0_dram_port_cmd_buffer_fifo_in_last, soc_hdmi_out0_dram_port_cmd_buffer_fifo_in_first, soc_hdmi_out0_dram_port_cmd_buffer_fifo_in_payload_sel};
assign {soc_hdmi_out0_dram_port_cmd_buffer_fifo_out_last, soc_hdmi_out0_dram_port_cmd_buffer_fifo_out_first, soc_hdmi_out0_dram_port_cmd_buffer_fifo_out_payload_sel} = soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_dout;
assign soc_hdmi_out0_dram_port_cmd_buffer_sink_ready = soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_writable;
assign soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_we = soc_hdmi_out0_dram_port_cmd_buffer_sink_valid;
assign soc_hdmi_out0_dram_port_cmd_buffer_fifo_in_first = soc_hdmi_out0_dram_port_cmd_buffer_sink_first;
assign soc_hdmi_out0_dram_port_cmd_buffer_fifo_in_last = soc_hdmi_out0_dram_port_cmd_buffer_sink_last;
assign soc_hdmi_out0_dram_port_cmd_buffer_fifo_in_payload_sel = soc_hdmi_out0_dram_port_cmd_buffer_sink_payload_sel;
assign soc_hdmi_out0_dram_port_cmd_buffer_source_valid = soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_readable;
assign soc_hdmi_out0_dram_port_cmd_buffer_source_first = soc_hdmi_out0_dram_port_cmd_buffer_fifo_out_first;
assign soc_hdmi_out0_dram_port_cmd_buffer_source_last = soc_hdmi_out0_dram_port_cmd_buffer_fifo_out_last;
assign soc_hdmi_out0_dram_port_cmd_buffer_source_payload_sel = soc_hdmi_out0_dram_port_cmd_buffer_fifo_out_payload_sel;
assign soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_re = soc_hdmi_out0_dram_port_cmd_buffer_source_ready;
always @(*) begin
	soc_hdmi_out0_dram_port_cmd_buffer_wrport_adr <= 2'd0;
	if (soc_hdmi_out0_dram_port_cmd_buffer_replace) begin
		soc_hdmi_out0_dram_port_cmd_buffer_wrport_adr <= (soc_hdmi_out0_dram_port_cmd_buffer_produce - 1'd1);
	end else begin
		soc_hdmi_out0_dram_port_cmd_buffer_wrport_adr <= soc_hdmi_out0_dram_port_cmd_buffer_produce;
	end
end
assign soc_hdmi_out0_dram_port_cmd_buffer_wrport_dat_w = soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_din;
assign soc_hdmi_out0_dram_port_cmd_buffer_wrport_we = (soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_we & (soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_writable | soc_hdmi_out0_dram_port_cmd_buffer_replace));
assign soc_hdmi_out0_dram_port_cmd_buffer_do_read = (soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_readable & soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_re);
assign soc_hdmi_out0_dram_port_cmd_buffer_rdport_adr = soc_hdmi_out0_dram_port_cmd_buffer_consume;
assign soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_dout = soc_hdmi_out0_dram_port_cmd_buffer_rdport_dat_r;
assign soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_writable = (soc_hdmi_out0_dram_port_cmd_buffer_level != 3'd4);
assign soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_readable = (soc_hdmi_out0_dram_port_cmd_buffer_level != 1'd0);
assign soc_hdmi_out0_dram_port_rdata_buffer_pipe_ce = (soc_hdmi_out0_dram_port_rdata_buffer_source_ready | (~soc_hdmi_out0_dram_port_rdata_buffer_valid_n));
assign soc_hdmi_out0_dram_port_rdata_buffer_sink_ready = soc_hdmi_out0_dram_port_rdata_buffer_pipe_ce;
assign soc_hdmi_out0_dram_port_rdata_buffer_source_valid = soc_hdmi_out0_dram_port_rdata_buffer_valid_n;
assign soc_hdmi_out0_dram_port_rdata_buffer_busy = (1'd0 | soc_hdmi_out0_dram_port_rdata_buffer_valid_n);
assign soc_hdmi_out0_dram_port_rdata_buffer_source_first = soc_hdmi_out0_dram_port_rdata_buffer_first_n;
assign soc_hdmi_out0_dram_port_rdata_buffer_source_last = soc_hdmi_out0_dram_port_rdata_buffer_last_n;
assign soc_hdmi_out0_dram_port_rdata_converter_converter_sink_valid = soc_hdmi_out0_dram_port_rdata_converter_sink_valid;
assign soc_hdmi_out0_dram_port_rdata_converter_converter_sink_first = soc_hdmi_out0_dram_port_rdata_converter_sink_first;
assign soc_hdmi_out0_dram_port_rdata_converter_converter_sink_last = soc_hdmi_out0_dram_port_rdata_converter_sink_last;
assign soc_hdmi_out0_dram_port_rdata_converter_sink_ready = soc_hdmi_out0_dram_port_rdata_converter_converter_sink_ready;
always @(*) begin
	soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data <= 128'd0;
	soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[15:0] <= soc_hdmi_out0_dram_port_rdata_converter_sink_payload_data[15:0];
	soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[31:16] <= soc_hdmi_out0_dram_port_rdata_converter_sink_payload_data[31:16];
	soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[47:32] <= soc_hdmi_out0_dram_port_rdata_converter_sink_payload_data[47:32];
	soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[63:48] <= soc_hdmi_out0_dram_port_rdata_converter_sink_payload_data[63:48];
	soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[79:64] <= soc_hdmi_out0_dram_port_rdata_converter_sink_payload_data[79:64];
	soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[95:80] <= soc_hdmi_out0_dram_port_rdata_converter_sink_payload_data[95:80];
	soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[111:96] <= soc_hdmi_out0_dram_port_rdata_converter_sink_payload_data[111:96];
	soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[127:112] <= soc_hdmi_out0_dram_port_rdata_converter_sink_payload_data[127:112];
end
assign soc_hdmi_out0_dram_port_rdata_converter_source_valid = soc_hdmi_out0_dram_port_rdata_converter_source_source_valid;
assign soc_hdmi_out0_dram_port_rdata_converter_source_first = soc_hdmi_out0_dram_port_rdata_converter_source_source_first;
assign soc_hdmi_out0_dram_port_rdata_converter_source_last = soc_hdmi_out0_dram_port_rdata_converter_source_source_last;
assign soc_hdmi_out0_dram_port_rdata_converter_source_source_ready = soc_hdmi_out0_dram_port_rdata_converter_source_ready;
assign {soc_hdmi_out0_dram_port_rdata_converter_source_payload_data} = soc_hdmi_out0_dram_port_rdata_converter_source_source_payload_data;
assign soc_hdmi_out0_dram_port_rdata_converter_source_source_valid = soc_hdmi_out0_dram_port_rdata_converter_converter_source_valid;
assign soc_hdmi_out0_dram_port_rdata_converter_converter_source_ready = soc_hdmi_out0_dram_port_rdata_converter_source_source_ready;
assign soc_hdmi_out0_dram_port_rdata_converter_source_source_first = soc_hdmi_out0_dram_port_rdata_converter_converter_source_first;
assign soc_hdmi_out0_dram_port_rdata_converter_source_source_last = soc_hdmi_out0_dram_port_rdata_converter_converter_source_last;
assign soc_hdmi_out0_dram_port_rdata_converter_source_source_payload_data = soc_hdmi_out0_dram_port_rdata_converter_converter_source_payload_data;
assign soc_hdmi_out0_dram_port_rdata_converter_converter_first = (soc_hdmi_out0_dram_port_rdata_converter_converter_mux == 1'd0);
assign soc_hdmi_out0_dram_port_rdata_converter_converter_last = (soc_hdmi_out0_dram_port_rdata_converter_converter_mux == 3'd7);
assign soc_hdmi_out0_dram_port_rdata_converter_converter_source_valid = soc_hdmi_out0_dram_port_rdata_converter_converter_sink_valid;
assign soc_hdmi_out0_dram_port_rdata_converter_converter_source_first = (soc_hdmi_out0_dram_port_rdata_converter_converter_sink_first & soc_hdmi_out0_dram_port_rdata_converter_converter_first);
assign soc_hdmi_out0_dram_port_rdata_converter_converter_source_last = (soc_hdmi_out0_dram_port_rdata_converter_converter_sink_last & soc_hdmi_out0_dram_port_rdata_converter_converter_last);
assign soc_hdmi_out0_dram_port_rdata_converter_converter_sink_ready = (soc_hdmi_out0_dram_port_rdata_converter_converter_last & soc_hdmi_out0_dram_port_rdata_converter_converter_source_ready);
always @(*) begin
	soc_hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= 16'd0;
	case (soc_hdmi_out0_dram_port_rdata_converter_converter_mux)
		1'd0: begin
			soc_hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[127:112];
		end
		1'd1: begin
			soc_hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[111:96];
		end
		2'd2: begin
			soc_hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[95:80];
		end
		2'd3: begin
			soc_hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[79:64];
		end
		3'd4: begin
			soc_hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[63:48];
		end
		3'd5: begin
			soc_hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[47:32];
		end
		3'd6: begin
			soc_hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[31:16];
		end
		default: begin
			soc_hdmi_out0_dram_port_rdata_converter_converter_source_payload_data <= soc_hdmi_out0_dram_port_rdata_converter_converter_sink_payload_data[15:0];
		end
	endcase
end
assign soc_hdmi_out0_dram_port_rdata_converter_converter_source_payload_valid_token_count = soc_hdmi_out0_dram_port_rdata_converter_converter_last;
assign soc_videosoc_data_port_adr = soc_videosoc_interface0_wb_sdram_adr[10:2];
always @(*) begin
	soc_videosoc_data_port_dat_w <= 128'd0;
	soc_videosoc_data_port_we <= 16'd0;
	if (soc_videosoc_write_from_slave) begin
		soc_videosoc_data_port_dat_w <= soc_videosoc_interface_dat_r;
		soc_videosoc_data_port_we <= {16{1'd1}};
	end else begin
		soc_videosoc_data_port_dat_w <= {4{soc_videosoc_interface0_wb_sdram_dat_w}};
		if ((((soc_videosoc_interface0_wb_sdram_cyc & soc_videosoc_interface0_wb_sdram_stb) & soc_videosoc_interface0_wb_sdram_we) & soc_videosoc_interface0_wb_sdram_ack)) begin
			soc_videosoc_data_port_we <= {({4{(soc_videosoc_interface0_wb_sdram_adr[1:0] == 1'd0)}} & soc_videosoc_interface0_wb_sdram_sel), ({4{(soc_videosoc_interface0_wb_sdram_adr[1:0] == 1'd1)}} & soc_videosoc_interface0_wb_sdram_sel), ({4{(soc_videosoc_interface0_wb_sdram_adr[1:0] == 2'd2)}} & soc_videosoc_interface0_wb_sdram_sel), ({4{(soc_videosoc_interface0_wb_sdram_adr[1:0] == 2'd3)}} & soc_videosoc_interface0_wb_sdram_sel)};
		end
	end
end
assign soc_videosoc_interface_dat_w = soc_videosoc_data_port_dat_r;
assign soc_videosoc_interface_sel = 16'd65535;
always @(*) begin
	soc_videosoc_interface0_wb_sdram_dat_r <= 32'd0;
	case (soc_videosoc_adr_offset_r)
		1'd0: begin
			soc_videosoc_interface0_wb_sdram_dat_r <= soc_videosoc_data_port_dat_r[127:96];
		end
		1'd1: begin
			soc_videosoc_interface0_wb_sdram_dat_r <= soc_videosoc_data_port_dat_r[95:64];
		end
		2'd2: begin
			soc_videosoc_interface0_wb_sdram_dat_r <= soc_videosoc_data_port_dat_r[63:32];
		end
		default: begin
			soc_videosoc_interface0_wb_sdram_dat_r <= soc_videosoc_data_port_dat_r[31:0];
		end
	endcase
end
assign {soc_videosoc_tag_do_dirty, soc_videosoc_tag_do_tag} = soc_videosoc_tag_port_dat_r;
assign soc_videosoc_tag_port_dat_w = {soc_videosoc_tag_di_dirty, soc_videosoc_tag_di_tag};
assign soc_videosoc_tag_port_adr = soc_videosoc_interface0_wb_sdram_adr[10:2];
assign soc_videosoc_tag_di_tag = soc_videosoc_interface0_wb_sdram_adr[29:11];
assign soc_videosoc_interface_adr = {soc_videosoc_tag_do_tag, soc_videosoc_interface0_wb_sdram_adr[10:2]};
always @(*) begin
	soc_videosoc_word_inc <= 1'd0;
	soc_videosoc_write_from_slave <= 1'd0;
	soc_videosoc_interface_cyc <= 1'd0;
	soc_videosoc_interface_stb <= 1'd0;
	soc_videosoc_tag_port_we <= 1'd0;
	soc_videosoc_interface0_wb_sdram_ack <= 1'd0;
	soc_videosoc_interface_we <= 1'd0;
	vns_fullmemorywe_next_state <= 3'd0;
	soc_videosoc_tag_di_dirty <= 1'd0;
	soc_videosoc_word_clr <= 1'd0;
	vns_fullmemorywe_next_state <= vns_fullmemorywe_state;
	case (vns_fullmemorywe_state)
		1'd1: begin
			soc_videosoc_word_clr <= 1'd1;
			if ((soc_videosoc_tag_do_tag == soc_videosoc_interface0_wb_sdram_adr[29:11])) begin
				soc_videosoc_interface0_wb_sdram_ack <= 1'd1;
				if (soc_videosoc_interface0_wb_sdram_we) begin
					soc_videosoc_tag_di_dirty <= 1'd1;
					soc_videosoc_tag_port_we <= 1'd1;
				end
				vns_fullmemorywe_next_state <= 1'd0;
			end else begin
				if (soc_videosoc_tag_do_dirty) begin
					vns_fullmemorywe_next_state <= 2'd2;
				end else begin
					vns_fullmemorywe_next_state <= 2'd3;
				end
			end
		end
		2'd2: begin
			soc_videosoc_interface_stb <= 1'd1;
			soc_videosoc_interface_cyc <= 1'd1;
			soc_videosoc_interface_we <= 1'd1;
			if (soc_videosoc_interface_ack) begin
				soc_videosoc_word_inc <= 1'd1;
				if (1'd1) begin
					vns_fullmemorywe_next_state <= 2'd3;
				end
			end
		end
		2'd3: begin
			soc_videosoc_tag_port_we <= 1'd1;
			soc_videosoc_word_clr <= 1'd1;
			vns_fullmemorywe_next_state <= 3'd4;
		end
		3'd4: begin
			soc_videosoc_interface_stb <= 1'd1;
			soc_videosoc_interface_cyc <= 1'd1;
			soc_videosoc_interface_we <= 1'd0;
			if (soc_videosoc_interface_ack) begin
				soc_videosoc_write_from_slave <= 1'd1;
				soc_videosoc_word_inc <= 1'd1;
				if (1'd1) begin
					vns_fullmemorywe_next_state <= 1'd1;
				end else begin
					vns_fullmemorywe_next_state <= 3'd4;
				end
			end
		end
		default: begin
			if ((soc_videosoc_interface0_wb_sdram_cyc & soc_videosoc_interface0_wb_sdram_stb)) begin
				vns_fullmemorywe_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_videosoc_port_cmd_payload_adr = soc_videosoc_interface_adr;
assign soc_videosoc_port_wdata_payload_we = soc_videosoc_interface_sel;
assign soc_videosoc_port_wdata_payload_data = soc_videosoc_interface_dat_w;
assign soc_videosoc_interface_dat_r = soc_videosoc_port_rdata_payload_data;
always @(*) begin
	soc_videosoc_port_cmd_payload_we <= 1'd0;
	soc_videosoc_port_rdata_ready <= 1'd0;
	vns_litedramwishbonebridge_next_state <= 2'd0;
	soc_videosoc_port_wdata_valid <= 1'd0;
	soc_videosoc_interface_ack <= 1'd0;
	soc_videosoc_port_cmd_valid <= 1'd0;
	vns_litedramwishbonebridge_next_state <= vns_litedramwishbonebridge_state;
	case (vns_litedramwishbonebridge_state)
		1'd1: begin
			soc_videosoc_port_cmd_valid <= 1'd1;
			soc_videosoc_port_cmd_payload_we <= soc_videosoc_interface_we;
			if (soc_videosoc_port_cmd_ready) begin
				if (soc_videosoc_interface_we) begin
					vns_litedramwishbonebridge_next_state <= 2'd2;
				end else begin
					vns_litedramwishbonebridge_next_state <= 2'd3;
				end
			end
		end
		2'd2: begin
			soc_videosoc_port_wdata_valid <= 1'd1;
			if (soc_videosoc_port_wdata_ready) begin
				soc_videosoc_interface_ack <= 1'd1;
				vns_litedramwishbonebridge_next_state <= 1'd0;
			end
		end
		2'd3: begin
			soc_videosoc_port_rdata_ready <= 1'd1;
			if (soc_videosoc_port_rdata_valid) begin
				soc_videosoc_interface_ack <= 1'd1;
				vns_litedramwishbonebridge_next_state <= 1'd0;
			end
		end
		default: begin
			if ((soc_videosoc_interface_cyc & soc_videosoc_interface_stb)) begin
				vns_litedramwishbonebridge_next_state <= 1'd1;
			end
		end
	endcase
end
assign spiflash_1x_wp = 1'd1;
assign spiflash_1x_hold = 1'd1;
assign soc_videosoc_bus_dat_r = soc_videosoc_sr;
always @(*) begin
	spiflash_1x_mosi <= 1'd0;
	spiflash_1x_cs_n <= 1'd0;
	soc_videosoc_clk0 <= 1'd0;
	soc_videosoc_miso_status <= 1'd0;
	if (soc_videosoc_bitbang_en_storage) begin
		soc_videosoc_clk0 <= soc_videosoc_bitbang_storage[1];
		spiflash_1x_cs_n <= soc_videosoc_bitbang_storage[2];
		if (soc_videosoc_bitbang_storage[1]) begin
			soc_videosoc_miso_status <= spiflash_1x_miso;
		end
		spiflash_1x_mosi <= soc_videosoc_bitbang_storage[0];
	end else begin
		soc_videosoc_clk0 <= soc_videosoc_clk1;
		spiflash_1x_cs_n <= soc_videosoc_cs_n;
		spiflash_1x_mosi <= soc_videosoc_sr[31];
	end
end
assign soc_ethphy_reset0 = (soc_ethphy_reset_storage | soc_ethphy_reset1);
assign eth_rst_n = (~soc_ethphy_reset0);
assign soc_ethphy_counter_done = (soc_ethphy_counter == 9'd256);
assign soc_ethphy_counter_ce = (~soc_ethphy_counter_done);
assign soc_ethphy_reset1 = (~soc_ethphy_counter_done);
assign soc_ethphy_sink_ready = 1'd1;
assign soc_ethphy_last = ((~soc_ethphy_rx_ctl) & soc_ethphy_rx_ctl_d);
assign soc_ethphy_source_last = soc_ethphy_last;
assign eth_mdc = soc_ethphy_storage[0];
assign soc_ethphy_data_oe = soc_ethphy_storage[1];
assign soc_ethphy_data_w = soc_ethphy_storage[2];
assign soc_ethmac_tx_cdc_sink_valid = soc_ethmac_source_valid;
assign soc_ethmac_source_ready = soc_ethmac_tx_cdc_sink_ready;
assign soc_ethmac_tx_cdc_sink_first = soc_ethmac_source_first;
assign soc_ethmac_tx_cdc_sink_last = soc_ethmac_source_last;
assign soc_ethmac_tx_cdc_sink_payload_data = soc_ethmac_source_payload_data;
assign soc_ethmac_tx_cdc_sink_payload_last_be = soc_ethmac_source_payload_last_be;
assign soc_ethmac_tx_cdc_sink_payload_error = soc_ethmac_source_payload_error;
assign soc_ethmac_sink_valid = soc_ethmac_rx_cdc_source_valid;
assign soc_ethmac_rx_cdc_source_ready = soc_ethmac_sink_ready;
assign soc_ethmac_sink_first = soc_ethmac_rx_cdc_source_first;
assign soc_ethmac_sink_last = soc_ethmac_rx_cdc_source_last;
assign soc_ethmac_sink_payload_data = soc_ethmac_rx_cdc_source_payload_data;
assign soc_ethmac_sink_payload_last_be = soc_ethmac_rx_cdc_source_payload_last_be;
assign soc_ethmac_sink_payload_error = soc_ethmac_rx_cdc_source_payload_error;
always @(*) begin
	soc_ethmac_tx_gap_inserter_source_payload_error <= 1'd0;
	soc_ethmac_tx_gap_inserter_counter_reset <= 1'd0;
	soc_ethmac_tx_gap_inserter_counter_ce <= 1'd0;
	soc_ethmac_tx_gap_inserter_sink_ready <= 1'd0;
	soc_ethmac_tx_gap_inserter_source_valid <= 1'd0;
	soc_ethmac_tx_gap_inserter_source_first <= 1'd0;
	vns_clockdomainsrenamer0_next_state <= 1'd0;
	soc_ethmac_tx_gap_inserter_source_last <= 1'd0;
	soc_ethmac_tx_gap_inserter_source_payload_data <= 8'd0;
	soc_ethmac_tx_gap_inserter_source_payload_last_be <= 1'd0;
	vns_clockdomainsrenamer0_next_state <= vns_clockdomainsrenamer0_state;
	case (vns_clockdomainsrenamer0_state)
		1'd1: begin
			soc_ethmac_tx_gap_inserter_counter_ce <= 1'd1;
			soc_ethmac_tx_gap_inserter_sink_ready <= 1'd0;
			if ((soc_ethmac_tx_gap_inserter_counter == 4'd11)) begin
				vns_clockdomainsrenamer0_next_state <= 1'd0;
			end
		end
		default: begin
			soc_ethmac_tx_gap_inserter_counter_reset <= 1'd1;
			soc_ethmac_tx_gap_inserter_source_valid <= soc_ethmac_tx_gap_inserter_sink_valid;
			soc_ethmac_tx_gap_inserter_sink_ready <= soc_ethmac_tx_gap_inserter_source_ready;
			soc_ethmac_tx_gap_inserter_source_first <= soc_ethmac_tx_gap_inserter_sink_first;
			soc_ethmac_tx_gap_inserter_source_last <= soc_ethmac_tx_gap_inserter_sink_last;
			soc_ethmac_tx_gap_inserter_source_payload_data <= soc_ethmac_tx_gap_inserter_sink_payload_data;
			soc_ethmac_tx_gap_inserter_source_payload_last_be <= soc_ethmac_tx_gap_inserter_sink_payload_last_be;
			soc_ethmac_tx_gap_inserter_source_payload_error <= soc_ethmac_tx_gap_inserter_sink_payload_error;
			if (((soc_ethmac_tx_gap_inserter_sink_valid & soc_ethmac_tx_gap_inserter_sink_last) & soc_ethmac_tx_gap_inserter_sink_ready)) begin
				vns_clockdomainsrenamer0_next_state <= 1'd1;
			end
		end
	endcase
end
always @(*) begin
	soc_ethmac_rx_gap_checker_source_valid <= 1'd0;
	soc_ethmac_rx_gap_checker_source_first <= 1'd0;
	soc_ethmac_rx_gap_checker_source_last <= 1'd0;
	vns_clockdomainsrenamer1_next_state <= 1'd0;
	soc_ethmac_rx_gap_checker_source_payload_data <= 8'd0;
	soc_ethmac_rx_gap_checker_source_payload_last_be <= 1'd0;
	soc_ethmac_rx_gap_checker_source_payload_error <= 1'd0;
	soc_ethmac_rx_gap_checker_counter_reset <= 1'd0;
	soc_ethmac_rx_gap_checker_counter_ce <= 1'd0;
	soc_ethmac_rx_gap_checker_sink_ready <= 1'd0;
	vns_clockdomainsrenamer1_next_state <= vns_clockdomainsrenamer1_state;
	case (vns_clockdomainsrenamer1_state)
		1'd1: begin
			soc_ethmac_rx_gap_checker_counter_ce <= 1'd1;
			soc_ethmac_rx_gap_checker_sink_ready <= 1'd1;
			if ((soc_ethmac_rx_gap_checker_counter == 4'd11)) begin
				vns_clockdomainsrenamer1_next_state <= 1'd0;
			end
		end
		default: begin
			soc_ethmac_rx_gap_checker_counter_reset <= 1'd1;
			soc_ethmac_rx_gap_checker_source_valid <= soc_ethmac_rx_gap_checker_sink_valid;
			soc_ethmac_rx_gap_checker_sink_ready <= soc_ethmac_rx_gap_checker_source_ready;
			soc_ethmac_rx_gap_checker_source_first <= soc_ethmac_rx_gap_checker_sink_first;
			soc_ethmac_rx_gap_checker_source_last <= soc_ethmac_rx_gap_checker_sink_last;
			soc_ethmac_rx_gap_checker_source_payload_data <= soc_ethmac_rx_gap_checker_sink_payload_data;
			soc_ethmac_rx_gap_checker_source_payload_last_be <= soc_ethmac_rx_gap_checker_sink_payload_last_be;
			soc_ethmac_rx_gap_checker_source_payload_error <= soc_ethmac_rx_gap_checker_sink_payload_error;
			if (((soc_ethmac_rx_gap_checker_sink_valid & soc_ethmac_rx_gap_checker_sink_last) & soc_ethmac_rx_gap_checker_sink_ready)) begin
				vns_clockdomainsrenamer1_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_ethmac_preamble_inserter_source_payload_last_be = soc_ethmac_preamble_inserter_sink_payload_last_be;
always @(*) begin
	soc_ethmac_preamble_inserter_clr_cnt <= 1'd0;
	soc_ethmac_preamble_inserter_inc_cnt <= 1'd0;
	soc_ethmac_preamble_inserter_sink_ready <= 1'd0;
	soc_ethmac_preamble_inserter_source_valid <= 1'd0;
	soc_ethmac_preamble_inserter_source_first <= 1'd0;
	vns_clockdomainsrenamer2_next_state <= 2'd0;
	soc_ethmac_preamble_inserter_source_last <= 1'd0;
	soc_ethmac_preamble_inserter_source_payload_data <= 8'd0;
	soc_ethmac_preamble_inserter_source_payload_error <= 1'd0;
	soc_ethmac_preamble_inserter_source_payload_data <= soc_ethmac_preamble_inserter_sink_payload_data;
	vns_clockdomainsrenamer2_next_state <= vns_clockdomainsrenamer2_state;
	case (vns_clockdomainsrenamer2_state)
		1'd1: begin
			soc_ethmac_preamble_inserter_source_valid <= 1'd1;
			case (soc_ethmac_preamble_inserter_cnt)
				1'd0: begin
					soc_ethmac_preamble_inserter_source_payload_data <= soc_ethmac_preamble_inserter_preamble[7:0];
				end
				1'd1: begin
					soc_ethmac_preamble_inserter_source_payload_data <= soc_ethmac_preamble_inserter_preamble[15:8];
				end
				2'd2: begin
					soc_ethmac_preamble_inserter_source_payload_data <= soc_ethmac_preamble_inserter_preamble[23:16];
				end
				2'd3: begin
					soc_ethmac_preamble_inserter_source_payload_data <= soc_ethmac_preamble_inserter_preamble[31:24];
				end
				3'd4: begin
					soc_ethmac_preamble_inserter_source_payload_data <= soc_ethmac_preamble_inserter_preamble[39:32];
				end
				3'd5: begin
					soc_ethmac_preamble_inserter_source_payload_data <= soc_ethmac_preamble_inserter_preamble[47:40];
				end
				3'd6: begin
					soc_ethmac_preamble_inserter_source_payload_data <= soc_ethmac_preamble_inserter_preamble[55:48];
				end
				default: begin
					soc_ethmac_preamble_inserter_source_payload_data <= soc_ethmac_preamble_inserter_preamble[63:56];
				end
			endcase
			if ((soc_ethmac_preamble_inserter_cnt == 3'd7)) begin
				if (soc_ethmac_preamble_inserter_source_ready) begin
					vns_clockdomainsrenamer2_next_state <= 2'd2;
				end
			end else begin
				soc_ethmac_preamble_inserter_inc_cnt <= soc_ethmac_preamble_inserter_source_ready;
			end
		end
		2'd2: begin
			soc_ethmac_preamble_inserter_source_valid <= soc_ethmac_preamble_inserter_sink_valid;
			soc_ethmac_preamble_inserter_sink_ready <= soc_ethmac_preamble_inserter_source_ready;
			soc_ethmac_preamble_inserter_source_first <= soc_ethmac_preamble_inserter_sink_first;
			soc_ethmac_preamble_inserter_source_last <= soc_ethmac_preamble_inserter_sink_last;
			soc_ethmac_preamble_inserter_source_payload_error <= soc_ethmac_preamble_inserter_sink_payload_error;
			if (((soc_ethmac_preamble_inserter_sink_valid & soc_ethmac_preamble_inserter_sink_last) & soc_ethmac_preamble_inserter_source_ready)) begin
				vns_clockdomainsrenamer2_next_state <= 1'd0;
			end
		end
		default: begin
			soc_ethmac_preamble_inserter_sink_ready <= 1'd1;
			soc_ethmac_preamble_inserter_clr_cnt <= 1'd1;
			if (soc_ethmac_preamble_inserter_sink_valid) begin
				soc_ethmac_preamble_inserter_sink_ready <= 1'd0;
				vns_clockdomainsrenamer2_next_state <= 1'd1;
			end
		end
	endcase
end
always @(*) begin
	soc_ethmac_preamble_checker_ref <= 8'd0;
	case (soc_ethmac_preamble_checker_cnt)
		1'd0: begin
			soc_ethmac_preamble_checker_ref <= soc_ethmac_preamble_checker_preamble[7:0];
		end
		1'd1: begin
			soc_ethmac_preamble_checker_ref <= soc_ethmac_preamble_checker_preamble[15:8];
		end
		2'd2: begin
			soc_ethmac_preamble_checker_ref <= soc_ethmac_preamble_checker_preamble[23:16];
		end
		2'd3: begin
			soc_ethmac_preamble_checker_ref <= soc_ethmac_preamble_checker_preamble[31:24];
		end
		3'd4: begin
			soc_ethmac_preamble_checker_ref <= soc_ethmac_preamble_checker_preamble[39:32];
		end
		3'd5: begin
			soc_ethmac_preamble_checker_ref <= soc_ethmac_preamble_checker_preamble[47:40];
		end
		3'd6: begin
			soc_ethmac_preamble_checker_ref <= soc_ethmac_preamble_checker_preamble[55:48];
		end
		default: begin
			soc_ethmac_preamble_checker_ref <= soc_ethmac_preamble_checker_preamble[63:56];
		end
	endcase
end
assign soc_ethmac_preamble_checker_match = (soc_ethmac_preamble_checker_sink_payload_data == soc_ethmac_preamble_checker_ref);
assign soc_ethmac_preamble_checker_source_payload_data = soc_ethmac_preamble_checker_sink_payload_data;
assign soc_ethmac_preamble_checker_source_payload_last_be = soc_ethmac_preamble_checker_sink_payload_last_be;
always @(*) begin
	soc_ethmac_preamble_checker_clr_cnt <= 1'd0;
	soc_ethmac_preamble_checker_sink_ready <= 1'd0;
	soc_ethmac_preamble_checker_inc_cnt <= 1'd0;
	soc_ethmac_preamble_checker_clr_discard <= 1'd0;
	soc_ethmac_preamble_checker_set_discard <= 1'd0;
	vns_clockdomainsrenamer3_next_state <= 2'd0;
	soc_ethmac_preamble_checker_source_valid <= 1'd0;
	soc_ethmac_preamble_checker_source_first <= 1'd0;
	soc_ethmac_preamble_checker_source_last <= 1'd0;
	soc_ethmac_preamble_checker_source_payload_error <= 1'd0;
	vns_clockdomainsrenamer3_next_state <= vns_clockdomainsrenamer3_state;
	case (vns_clockdomainsrenamer3_state)
		1'd1: begin
			soc_ethmac_preamble_checker_sink_ready <= 1'd1;
			if (soc_ethmac_preamble_checker_sink_valid) begin
				soc_ethmac_preamble_checker_set_discard <= (~soc_ethmac_preamble_checker_match);
				if ((soc_ethmac_preamble_checker_cnt == 3'd7)) begin
					if ((soc_ethmac_preamble_checker_discard | (~soc_ethmac_preamble_checker_match))) begin
						vns_clockdomainsrenamer3_next_state <= 1'd0;
					end else begin
						vns_clockdomainsrenamer3_next_state <= 2'd2;
					end
				end else begin
					soc_ethmac_preamble_checker_inc_cnt <= 1'd1;
				end
			end
		end
		2'd2: begin
			soc_ethmac_preamble_checker_source_valid <= soc_ethmac_preamble_checker_sink_valid;
			soc_ethmac_preamble_checker_sink_ready <= soc_ethmac_preamble_checker_source_ready;
			soc_ethmac_preamble_checker_source_first <= soc_ethmac_preamble_checker_sink_first;
			soc_ethmac_preamble_checker_source_last <= soc_ethmac_preamble_checker_sink_last;
			soc_ethmac_preamble_checker_source_payload_error <= soc_ethmac_preamble_checker_sink_payload_error;
			if (((soc_ethmac_preamble_checker_source_valid & soc_ethmac_preamble_checker_source_last) & soc_ethmac_preamble_checker_source_ready)) begin
				vns_clockdomainsrenamer3_next_state <= 1'd0;
			end
		end
		default: begin
			soc_ethmac_preamble_checker_sink_ready <= 1'd1;
			soc_ethmac_preamble_checker_clr_cnt <= 1'd1;
			soc_ethmac_preamble_checker_clr_discard <= 1'd1;
			if (soc_ethmac_preamble_checker_sink_valid) begin
				soc_ethmac_preamble_checker_clr_cnt <= 1'd0;
				soc_ethmac_preamble_checker_inc_cnt <= 1'd1;
				soc_ethmac_preamble_checker_clr_discard <= 1'd0;
				soc_ethmac_preamble_checker_set_discard <= (~soc_ethmac_preamble_checker_match);
				vns_clockdomainsrenamer3_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_ethmac_crc32_inserter_cnt_done = (soc_ethmac_crc32_inserter_cnt == 1'd0);
assign soc_ethmac_crc32_inserter_data1 = soc_ethmac_crc32_inserter_data0;
assign soc_ethmac_crc32_inserter_last = soc_ethmac_crc32_inserter_reg;
assign soc_ethmac_crc32_inserter_value = (~{soc_ethmac_crc32_inserter_reg[0], soc_ethmac_crc32_inserter_reg[1], soc_ethmac_crc32_inserter_reg[2], soc_ethmac_crc32_inserter_reg[3], soc_ethmac_crc32_inserter_reg[4], soc_ethmac_crc32_inserter_reg[5], soc_ethmac_crc32_inserter_reg[6], soc_ethmac_crc32_inserter_reg[7], soc_ethmac_crc32_inserter_reg[8], soc_ethmac_crc32_inserter_reg[9], soc_ethmac_crc32_inserter_reg[10], soc_ethmac_crc32_inserter_reg[11], soc_ethmac_crc32_inserter_reg[12], soc_ethmac_crc32_inserter_reg[13], soc_ethmac_crc32_inserter_reg[14], soc_ethmac_crc32_inserter_reg[15], soc_ethmac_crc32_inserter_reg[16], soc_ethmac_crc32_inserter_reg[17], soc_ethmac_crc32_inserter_reg[18], soc_ethmac_crc32_inserter_reg[19], soc_ethmac_crc32_inserter_reg[20], soc_ethmac_crc32_inserter_reg[21], soc_ethmac_crc32_inserter_reg[22], soc_ethmac_crc32_inserter_reg[23], soc_ethmac_crc32_inserter_reg[24], soc_ethmac_crc32_inserter_reg[25], soc_ethmac_crc32_inserter_reg[26], soc_ethmac_crc32_inserter_reg[27], soc_ethmac_crc32_inserter_reg[28], soc_ethmac_crc32_inserter_reg[29], soc_ethmac_crc32_inserter_reg[30], soc_ethmac_crc32_inserter_reg[31]});
assign soc_ethmac_crc32_inserter_error = (soc_ethmac_crc32_inserter_next != 32'd3338984827);
always @(*) begin
	soc_ethmac_crc32_inserter_next <= 32'd0;
	soc_ethmac_crc32_inserter_next[0] <= (((soc_ethmac_crc32_inserter_last[24] ^ soc_ethmac_crc32_inserter_last[30]) ^ soc_ethmac_crc32_inserter_data1[1]) ^ soc_ethmac_crc32_inserter_data1[7]);
	soc_ethmac_crc32_inserter_next[1] <= (((((((soc_ethmac_crc32_inserter_last[25] ^ soc_ethmac_crc32_inserter_last[31]) ^ soc_ethmac_crc32_inserter_data1[0]) ^ soc_ethmac_crc32_inserter_data1[6]) ^ soc_ethmac_crc32_inserter_last[24]) ^ soc_ethmac_crc32_inserter_last[30]) ^ soc_ethmac_crc32_inserter_data1[1]) ^ soc_ethmac_crc32_inserter_data1[7]);
	soc_ethmac_crc32_inserter_next[2] <= (((((((((soc_ethmac_crc32_inserter_last[26] ^ soc_ethmac_crc32_inserter_data1[5]) ^ soc_ethmac_crc32_inserter_last[25]) ^ soc_ethmac_crc32_inserter_last[31]) ^ soc_ethmac_crc32_inserter_data1[0]) ^ soc_ethmac_crc32_inserter_data1[6]) ^ soc_ethmac_crc32_inserter_last[24]) ^ soc_ethmac_crc32_inserter_last[30]) ^ soc_ethmac_crc32_inserter_data1[1]) ^ soc_ethmac_crc32_inserter_data1[7]);
	soc_ethmac_crc32_inserter_next[3] <= (((((((soc_ethmac_crc32_inserter_last[27] ^ soc_ethmac_crc32_inserter_data1[4]) ^ soc_ethmac_crc32_inserter_last[26]) ^ soc_ethmac_crc32_inserter_data1[5]) ^ soc_ethmac_crc32_inserter_last[25]) ^ soc_ethmac_crc32_inserter_last[31]) ^ soc_ethmac_crc32_inserter_data1[0]) ^ soc_ethmac_crc32_inserter_data1[6]);
	soc_ethmac_crc32_inserter_next[4] <= (((((((((soc_ethmac_crc32_inserter_last[28] ^ soc_ethmac_crc32_inserter_data1[3]) ^ soc_ethmac_crc32_inserter_last[27]) ^ soc_ethmac_crc32_inserter_data1[4]) ^ soc_ethmac_crc32_inserter_last[26]) ^ soc_ethmac_crc32_inserter_data1[5]) ^ soc_ethmac_crc32_inserter_last[24]) ^ soc_ethmac_crc32_inserter_last[30]) ^ soc_ethmac_crc32_inserter_data1[1]) ^ soc_ethmac_crc32_inserter_data1[7]);
	soc_ethmac_crc32_inserter_next[5] <= (((((((((((((soc_ethmac_crc32_inserter_last[29] ^ soc_ethmac_crc32_inserter_data1[2]) ^ soc_ethmac_crc32_inserter_last[28]) ^ soc_ethmac_crc32_inserter_data1[3]) ^ soc_ethmac_crc32_inserter_last[27]) ^ soc_ethmac_crc32_inserter_data1[4]) ^ soc_ethmac_crc32_inserter_last[25]) ^ soc_ethmac_crc32_inserter_last[31]) ^ soc_ethmac_crc32_inserter_data1[0]) ^ soc_ethmac_crc32_inserter_data1[6]) ^ soc_ethmac_crc32_inserter_last[24]) ^ soc_ethmac_crc32_inserter_last[30]) ^ soc_ethmac_crc32_inserter_data1[1]) ^ soc_ethmac_crc32_inserter_data1[7]);
	soc_ethmac_crc32_inserter_next[6] <= (((((((((((soc_ethmac_crc32_inserter_last[30] ^ soc_ethmac_crc32_inserter_data1[1]) ^ soc_ethmac_crc32_inserter_last[29]) ^ soc_ethmac_crc32_inserter_data1[2]) ^ soc_ethmac_crc32_inserter_last[28]) ^ soc_ethmac_crc32_inserter_data1[3]) ^ soc_ethmac_crc32_inserter_last[26]) ^ soc_ethmac_crc32_inserter_data1[5]) ^ soc_ethmac_crc32_inserter_last[25]) ^ soc_ethmac_crc32_inserter_last[31]) ^ soc_ethmac_crc32_inserter_data1[0]) ^ soc_ethmac_crc32_inserter_data1[6]);
	soc_ethmac_crc32_inserter_next[7] <= (((((((((soc_ethmac_crc32_inserter_last[31] ^ soc_ethmac_crc32_inserter_data1[0]) ^ soc_ethmac_crc32_inserter_last[29]) ^ soc_ethmac_crc32_inserter_data1[2]) ^ soc_ethmac_crc32_inserter_last[27]) ^ soc_ethmac_crc32_inserter_data1[4]) ^ soc_ethmac_crc32_inserter_last[26]) ^ soc_ethmac_crc32_inserter_data1[5]) ^ soc_ethmac_crc32_inserter_last[24]) ^ soc_ethmac_crc32_inserter_data1[7]);
	soc_ethmac_crc32_inserter_next[8] <= ((((((((soc_ethmac_crc32_inserter_last[0] ^ soc_ethmac_crc32_inserter_last[28]) ^ soc_ethmac_crc32_inserter_data1[3]) ^ soc_ethmac_crc32_inserter_last[27]) ^ soc_ethmac_crc32_inserter_data1[4]) ^ soc_ethmac_crc32_inserter_last[25]) ^ soc_ethmac_crc32_inserter_data1[6]) ^ soc_ethmac_crc32_inserter_last[24]) ^ soc_ethmac_crc32_inserter_data1[7]);
	soc_ethmac_crc32_inserter_next[9] <= ((((((((soc_ethmac_crc32_inserter_last[1] ^ soc_ethmac_crc32_inserter_last[29]) ^ soc_ethmac_crc32_inserter_data1[2]) ^ soc_ethmac_crc32_inserter_last[28]) ^ soc_ethmac_crc32_inserter_data1[3]) ^ soc_ethmac_crc32_inserter_last[26]) ^ soc_ethmac_crc32_inserter_data1[5]) ^ soc_ethmac_crc32_inserter_last[25]) ^ soc_ethmac_crc32_inserter_data1[6]);
	soc_ethmac_crc32_inserter_next[10] <= ((((((((soc_ethmac_crc32_inserter_last[2] ^ soc_ethmac_crc32_inserter_last[29]) ^ soc_ethmac_crc32_inserter_data1[2]) ^ soc_ethmac_crc32_inserter_last[27]) ^ soc_ethmac_crc32_inserter_data1[4]) ^ soc_ethmac_crc32_inserter_last[26]) ^ soc_ethmac_crc32_inserter_data1[5]) ^ soc_ethmac_crc32_inserter_last[24]) ^ soc_ethmac_crc32_inserter_data1[7]);
	soc_ethmac_crc32_inserter_next[11] <= ((((((((soc_ethmac_crc32_inserter_last[3] ^ soc_ethmac_crc32_inserter_last[28]) ^ soc_ethmac_crc32_inserter_data1[3]) ^ soc_ethmac_crc32_inserter_last[27]) ^ soc_ethmac_crc32_inserter_data1[4]) ^ soc_ethmac_crc32_inserter_last[25]) ^ soc_ethmac_crc32_inserter_data1[6]) ^ soc_ethmac_crc32_inserter_last[24]) ^ soc_ethmac_crc32_inserter_data1[7]);
	soc_ethmac_crc32_inserter_next[12] <= ((((((((((((soc_ethmac_crc32_inserter_last[4] ^ soc_ethmac_crc32_inserter_last[29]) ^ soc_ethmac_crc32_inserter_data1[2]) ^ soc_ethmac_crc32_inserter_last[28]) ^ soc_ethmac_crc32_inserter_data1[3]) ^ soc_ethmac_crc32_inserter_last[26]) ^ soc_ethmac_crc32_inserter_data1[5]) ^ soc_ethmac_crc32_inserter_last[25]) ^ soc_ethmac_crc32_inserter_data1[6]) ^ soc_ethmac_crc32_inserter_last[24]) ^ soc_ethmac_crc32_inserter_last[30]) ^ soc_ethmac_crc32_inserter_data1[1]) ^ soc_ethmac_crc32_inserter_data1[7]);
	soc_ethmac_crc32_inserter_next[13] <= ((((((((((((soc_ethmac_crc32_inserter_last[5] ^ soc_ethmac_crc32_inserter_last[30]) ^ soc_ethmac_crc32_inserter_data1[1]) ^ soc_ethmac_crc32_inserter_last[29]) ^ soc_ethmac_crc32_inserter_data1[2]) ^ soc_ethmac_crc32_inserter_last[27]) ^ soc_ethmac_crc32_inserter_data1[4]) ^ soc_ethmac_crc32_inserter_last[26]) ^ soc_ethmac_crc32_inserter_data1[5]) ^ soc_ethmac_crc32_inserter_last[25]) ^ soc_ethmac_crc32_inserter_last[31]) ^ soc_ethmac_crc32_inserter_data1[0]) ^ soc_ethmac_crc32_inserter_data1[6]);
	soc_ethmac_crc32_inserter_next[14] <= ((((((((((soc_ethmac_crc32_inserter_last[6] ^ soc_ethmac_crc32_inserter_last[31]) ^ soc_ethmac_crc32_inserter_data1[0]) ^ soc_ethmac_crc32_inserter_last[30]) ^ soc_ethmac_crc32_inserter_data1[1]) ^ soc_ethmac_crc32_inserter_last[28]) ^ soc_ethmac_crc32_inserter_data1[3]) ^ soc_ethmac_crc32_inserter_last[27]) ^ soc_ethmac_crc32_inserter_data1[4]) ^ soc_ethmac_crc32_inserter_last[26]) ^ soc_ethmac_crc32_inserter_data1[5]);
	soc_ethmac_crc32_inserter_next[15] <= ((((((((soc_ethmac_crc32_inserter_last[7] ^ soc_ethmac_crc32_inserter_last[31]) ^ soc_ethmac_crc32_inserter_data1[0]) ^ soc_ethmac_crc32_inserter_last[29]) ^ soc_ethmac_crc32_inserter_data1[2]) ^ soc_ethmac_crc32_inserter_last[28]) ^ soc_ethmac_crc32_inserter_data1[3]) ^ soc_ethmac_crc32_inserter_last[27]) ^ soc_ethmac_crc32_inserter_data1[4]);
	soc_ethmac_crc32_inserter_next[16] <= ((((((soc_ethmac_crc32_inserter_last[8] ^ soc_ethmac_crc32_inserter_last[29]) ^ soc_ethmac_crc32_inserter_data1[2]) ^ soc_ethmac_crc32_inserter_last[28]) ^ soc_ethmac_crc32_inserter_data1[3]) ^ soc_ethmac_crc32_inserter_last[24]) ^ soc_ethmac_crc32_inserter_data1[7]);
	soc_ethmac_crc32_inserter_next[17] <= ((((((soc_ethmac_crc32_inserter_last[9] ^ soc_ethmac_crc32_inserter_last[30]) ^ soc_ethmac_crc32_inserter_data1[1]) ^ soc_ethmac_crc32_inserter_last[29]) ^ soc_ethmac_crc32_inserter_data1[2]) ^ soc_ethmac_crc32_inserter_last[25]) ^ soc_ethmac_crc32_inserter_data1[6]);
	soc_ethmac_crc32_inserter_next[18] <= ((((((soc_ethmac_crc32_inserter_last[10] ^ soc_ethmac_crc32_inserter_last[31]) ^ soc_ethmac_crc32_inserter_data1[0]) ^ soc_ethmac_crc32_inserter_last[30]) ^ soc_ethmac_crc32_inserter_data1[1]) ^ soc_ethmac_crc32_inserter_last[26]) ^ soc_ethmac_crc32_inserter_data1[5]);
	soc_ethmac_crc32_inserter_next[19] <= ((((soc_ethmac_crc32_inserter_last[11] ^ soc_ethmac_crc32_inserter_last[31]) ^ soc_ethmac_crc32_inserter_data1[0]) ^ soc_ethmac_crc32_inserter_last[27]) ^ soc_ethmac_crc32_inserter_data1[4]);
	soc_ethmac_crc32_inserter_next[20] <= ((soc_ethmac_crc32_inserter_last[12] ^ soc_ethmac_crc32_inserter_last[28]) ^ soc_ethmac_crc32_inserter_data1[3]);
	soc_ethmac_crc32_inserter_next[21] <= ((soc_ethmac_crc32_inserter_last[13] ^ soc_ethmac_crc32_inserter_last[29]) ^ soc_ethmac_crc32_inserter_data1[2]);
	soc_ethmac_crc32_inserter_next[22] <= ((soc_ethmac_crc32_inserter_last[14] ^ soc_ethmac_crc32_inserter_last[24]) ^ soc_ethmac_crc32_inserter_data1[7]);
	soc_ethmac_crc32_inserter_next[23] <= ((((((soc_ethmac_crc32_inserter_last[15] ^ soc_ethmac_crc32_inserter_last[25]) ^ soc_ethmac_crc32_inserter_data1[6]) ^ soc_ethmac_crc32_inserter_last[24]) ^ soc_ethmac_crc32_inserter_last[30]) ^ soc_ethmac_crc32_inserter_data1[1]) ^ soc_ethmac_crc32_inserter_data1[7]);
	soc_ethmac_crc32_inserter_next[24] <= ((((((soc_ethmac_crc32_inserter_last[16] ^ soc_ethmac_crc32_inserter_last[26]) ^ soc_ethmac_crc32_inserter_data1[5]) ^ soc_ethmac_crc32_inserter_last[25]) ^ soc_ethmac_crc32_inserter_last[31]) ^ soc_ethmac_crc32_inserter_data1[0]) ^ soc_ethmac_crc32_inserter_data1[6]);
	soc_ethmac_crc32_inserter_next[25] <= ((((soc_ethmac_crc32_inserter_last[17] ^ soc_ethmac_crc32_inserter_last[27]) ^ soc_ethmac_crc32_inserter_data1[4]) ^ soc_ethmac_crc32_inserter_last[26]) ^ soc_ethmac_crc32_inserter_data1[5]);
	soc_ethmac_crc32_inserter_next[26] <= ((((((((soc_ethmac_crc32_inserter_last[18] ^ soc_ethmac_crc32_inserter_last[28]) ^ soc_ethmac_crc32_inserter_data1[3]) ^ soc_ethmac_crc32_inserter_last[27]) ^ soc_ethmac_crc32_inserter_data1[4]) ^ soc_ethmac_crc32_inserter_last[24]) ^ soc_ethmac_crc32_inserter_last[30]) ^ soc_ethmac_crc32_inserter_data1[1]) ^ soc_ethmac_crc32_inserter_data1[7]);
	soc_ethmac_crc32_inserter_next[27] <= ((((((((soc_ethmac_crc32_inserter_last[19] ^ soc_ethmac_crc32_inserter_last[29]) ^ soc_ethmac_crc32_inserter_data1[2]) ^ soc_ethmac_crc32_inserter_last[28]) ^ soc_ethmac_crc32_inserter_data1[3]) ^ soc_ethmac_crc32_inserter_last[25]) ^ soc_ethmac_crc32_inserter_last[31]) ^ soc_ethmac_crc32_inserter_data1[0]) ^ soc_ethmac_crc32_inserter_data1[6]);
	soc_ethmac_crc32_inserter_next[28] <= ((((((soc_ethmac_crc32_inserter_last[20] ^ soc_ethmac_crc32_inserter_last[30]) ^ soc_ethmac_crc32_inserter_data1[1]) ^ soc_ethmac_crc32_inserter_last[29]) ^ soc_ethmac_crc32_inserter_data1[2]) ^ soc_ethmac_crc32_inserter_last[26]) ^ soc_ethmac_crc32_inserter_data1[5]);
	soc_ethmac_crc32_inserter_next[29] <= ((((((soc_ethmac_crc32_inserter_last[21] ^ soc_ethmac_crc32_inserter_last[31]) ^ soc_ethmac_crc32_inserter_data1[0]) ^ soc_ethmac_crc32_inserter_last[30]) ^ soc_ethmac_crc32_inserter_data1[1]) ^ soc_ethmac_crc32_inserter_last[27]) ^ soc_ethmac_crc32_inserter_data1[4]);
	soc_ethmac_crc32_inserter_next[30] <= ((((soc_ethmac_crc32_inserter_last[22] ^ soc_ethmac_crc32_inserter_last[31]) ^ soc_ethmac_crc32_inserter_data1[0]) ^ soc_ethmac_crc32_inserter_last[28]) ^ soc_ethmac_crc32_inserter_data1[3]);
	soc_ethmac_crc32_inserter_next[31] <= ((soc_ethmac_crc32_inserter_last[23] ^ soc_ethmac_crc32_inserter_last[29]) ^ soc_ethmac_crc32_inserter_data1[2]);
end
always @(*) begin
	soc_ethmac_crc32_inserter_source_valid <= 1'd0;
	vns_clockdomainsrenamer4_next_state <= 2'd0;
	soc_ethmac_crc32_inserter_source_first <= 1'd0;
	soc_ethmac_crc32_inserter_source_last <= 1'd0;
	soc_ethmac_crc32_inserter_source_payload_data <= 8'd0;
	soc_ethmac_crc32_inserter_source_payload_last_be <= 1'd0;
	soc_ethmac_crc32_inserter_source_payload_error <= 1'd0;
	soc_ethmac_crc32_inserter_data0 <= 8'd0;
	soc_ethmac_crc32_inserter_is_ongoing0 <= 1'd0;
	soc_ethmac_crc32_inserter_sink_ready <= 1'd0;
	soc_ethmac_crc32_inserter_is_ongoing1 <= 1'd0;
	soc_ethmac_crc32_inserter_ce <= 1'd0;
	soc_ethmac_crc32_inserter_reset <= 1'd0;
	vns_clockdomainsrenamer4_next_state <= vns_clockdomainsrenamer4_state;
	case (vns_clockdomainsrenamer4_state)
		1'd1: begin
			soc_ethmac_crc32_inserter_ce <= (soc_ethmac_crc32_inserter_sink_valid & soc_ethmac_crc32_inserter_source_ready);
			soc_ethmac_crc32_inserter_data0 <= soc_ethmac_crc32_inserter_sink_payload_data;
			soc_ethmac_crc32_inserter_source_valid <= soc_ethmac_crc32_inserter_sink_valid;
			soc_ethmac_crc32_inserter_sink_ready <= soc_ethmac_crc32_inserter_source_ready;
			soc_ethmac_crc32_inserter_source_first <= soc_ethmac_crc32_inserter_sink_first;
			soc_ethmac_crc32_inserter_source_last <= soc_ethmac_crc32_inserter_sink_last;
			soc_ethmac_crc32_inserter_source_payload_data <= soc_ethmac_crc32_inserter_sink_payload_data;
			soc_ethmac_crc32_inserter_source_payload_last_be <= soc_ethmac_crc32_inserter_sink_payload_last_be;
			soc_ethmac_crc32_inserter_source_payload_error <= soc_ethmac_crc32_inserter_sink_payload_error;
			soc_ethmac_crc32_inserter_source_last <= 1'd0;
			if (((soc_ethmac_crc32_inserter_sink_valid & soc_ethmac_crc32_inserter_sink_last) & soc_ethmac_crc32_inserter_source_ready)) begin
				vns_clockdomainsrenamer4_next_state <= 2'd2;
			end
		end
		2'd2: begin
			soc_ethmac_crc32_inserter_source_valid <= 1'd1;
			case (soc_ethmac_crc32_inserter_cnt)
				1'd0: begin
					soc_ethmac_crc32_inserter_source_payload_data <= soc_ethmac_crc32_inserter_value[31:24];
				end
				1'd1: begin
					soc_ethmac_crc32_inserter_source_payload_data <= soc_ethmac_crc32_inserter_value[23:16];
				end
				2'd2: begin
					soc_ethmac_crc32_inserter_source_payload_data <= soc_ethmac_crc32_inserter_value[15:8];
				end
				default: begin
					soc_ethmac_crc32_inserter_source_payload_data <= soc_ethmac_crc32_inserter_value[7:0];
				end
			endcase
			if (soc_ethmac_crc32_inserter_cnt_done) begin
				soc_ethmac_crc32_inserter_source_last <= 1'd1;
				if (soc_ethmac_crc32_inserter_source_ready) begin
					vns_clockdomainsrenamer4_next_state <= 1'd0;
				end
			end
			soc_ethmac_crc32_inserter_is_ongoing1 <= 1'd1;
		end
		default: begin
			soc_ethmac_crc32_inserter_reset <= 1'd1;
			soc_ethmac_crc32_inserter_sink_ready <= 1'd1;
			if (soc_ethmac_crc32_inserter_sink_valid) begin
				soc_ethmac_crc32_inserter_sink_ready <= 1'd0;
				vns_clockdomainsrenamer4_next_state <= 1'd1;
			end
			soc_ethmac_crc32_inserter_is_ongoing0 <= 1'd1;
		end
	endcase
end
assign soc_ethmac_crc32_checker_fifo_full = (soc_ethmac_crc32_checker_syncfifo_level == 3'd4);
assign soc_ethmac_crc32_checker_fifo_in = (soc_ethmac_crc32_checker_sink_sink_valid & ((~soc_ethmac_crc32_checker_fifo_full) | soc_ethmac_crc32_checker_fifo_out));
assign soc_ethmac_crc32_checker_fifo_out = (soc_ethmac_crc32_checker_source_source_valid & soc_ethmac_crc32_checker_source_source_ready);
assign soc_ethmac_crc32_checker_syncfifo_sink_first = soc_ethmac_crc32_checker_sink_sink_first;
assign soc_ethmac_crc32_checker_syncfifo_sink_last = soc_ethmac_crc32_checker_sink_sink_last;
assign soc_ethmac_crc32_checker_syncfifo_sink_payload_data = soc_ethmac_crc32_checker_sink_sink_payload_data;
assign soc_ethmac_crc32_checker_syncfifo_sink_payload_last_be = soc_ethmac_crc32_checker_sink_sink_payload_last_be;
assign soc_ethmac_crc32_checker_syncfifo_sink_payload_error = soc_ethmac_crc32_checker_sink_sink_payload_error;
always @(*) begin
	soc_ethmac_crc32_checker_syncfifo_sink_valid <= 1'd0;
	soc_ethmac_crc32_checker_syncfifo_sink_valid <= soc_ethmac_crc32_checker_sink_sink_valid;
	soc_ethmac_crc32_checker_syncfifo_sink_valid <= soc_ethmac_crc32_checker_fifo_in;
end
always @(*) begin
	soc_ethmac_crc32_checker_sink_sink_ready <= 1'd0;
	soc_ethmac_crc32_checker_sink_sink_ready <= soc_ethmac_crc32_checker_syncfifo_sink_ready;
	soc_ethmac_crc32_checker_sink_sink_ready <= soc_ethmac_crc32_checker_fifo_in;
end
assign soc_ethmac_crc32_checker_source_source_valid = (soc_ethmac_crc32_checker_sink_sink_valid & soc_ethmac_crc32_checker_fifo_full);
assign soc_ethmac_crc32_checker_source_source_last = soc_ethmac_crc32_checker_sink_sink_last;
assign soc_ethmac_crc32_checker_syncfifo_source_ready = soc_ethmac_crc32_checker_fifo_out;
assign soc_ethmac_crc32_checker_source_source_payload_data = soc_ethmac_crc32_checker_syncfifo_source_payload_data;
assign soc_ethmac_crc32_checker_source_source_payload_last_be = soc_ethmac_crc32_checker_syncfifo_source_payload_last_be;
always @(*) begin
	soc_ethmac_crc32_checker_source_source_payload_error <= 1'd0;
	soc_ethmac_crc32_checker_source_source_payload_error <= soc_ethmac_crc32_checker_syncfifo_source_payload_error;
	soc_ethmac_crc32_checker_source_source_payload_error <= (soc_ethmac_crc32_checker_sink_sink_payload_error | soc_ethmac_crc32_checker_crc_error);
end
assign soc_ethmac_crc32_checker_crc_data0 = soc_ethmac_crc32_checker_sink_sink_payload_data;
assign soc_ethmac_crc32_checker_crc_data1 = soc_ethmac_crc32_checker_crc_data0;
assign soc_ethmac_crc32_checker_crc_last = soc_ethmac_crc32_checker_crc_reg;
assign soc_ethmac_crc32_checker_crc_value = (~{soc_ethmac_crc32_checker_crc_reg[0], soc_ethmac_crc32_checker_crc_reg[1], soc_ethmac_crc32_checker_crc_reg[2], soc_ethmac_crc32_checker_crc_reg[3], soc_ethmac_crc32_checker_crc_reg[4], soc_ethmac_crc32_checker_crc_reg[5], soc_ethmac_crc32_checker_crc_reg[6], soc_ethmac_crc32_checker_crc_reg[7], soc_ethmac_crc32_checker_crc_reg[8], soc_ethmac_crc32_checker_crc_reg[9], soc_ethmac_crc32_checker_crc_reg[10], soc_ethmac_crc32_checker_crc_reg[11], soc_ethmac_crc32_checker_crc_reg[12], soc_ethmac_crc32_checker_crc_reg[13], soc_ethmac_crc32_checker_crc_reg[14], soc_ethmac_crc32_checker_crc_reg[15], soc_ethmac_crc32_checker_crc_reg[16], soc_ethmac_crc32_checker_crc_reg[17], soc_ethmac_crc32_checker_crc_reg[18], soc_ethmac_crc32_checker_crc_reg[19], soc_ethmac_crc32_checker_crc_reg[20], soc_ethmac_crc32_checker_crc_reg[21], soc_ethmac_crc32_checker_crc_reg[22], soc_ethmac_crc32_checker_crc_reg[23], soc_ethmac_crc32_checker_crc_reg[24], soc_ethmac_crc32_checker_crc_reg[25], soc_ethmac_crc32_checker_crc_reg[26], soc_ethmac_crc32_checker_crc_reg[27], soc_ethmac_crc32_checker_crc_reg[28], soc_ethmac_crc32_checker_crc_reg[29], soc_ethmac_crc32_checker_crc_reg[30], soc_ethmac_crc32_checker_crc_reg[31]});
assign soc_ethmac_crc32_checker_crc_error = (soc_ethmac_crc32_checker_crc_next != 32'd3338984827);
always @(*) begin
	soc_ethmac_crc32_checker_crc_next <= 32'd0;
	soc_ethmac_crc32_checker_crc_next[0] <= (((soc_ethmac_crc32_checker_crc_last[24] ^ soc_ethmac_crc32_checker_crc_last[30]) ^ soc_ethmac_crc32_checker_crc_data1[1]) ^ soc_ethmac_crc32_checker_crc_data1[7]);
	soc_ethmac_crc32_checker_crc_next[1] <= (((((((soc_ethmac_crc32_checker_crc_last[25] ^ soc_ethmac_crc32_checker_crc_last[31]) ^ soc_ethmac_crc32_checker_crc_data1[0]) ^ soc_ethmac_crc32_checker_crc_data1[6]) ^ soc_ethmac_crc32_checker_crc_last[24]) ^ soc_ethmac_crc32_checker_crc_last[30]) ^ soc_ethmac_crc32_checker_crc_data1[1]) ^ soc_ethmac_crc32_checker_crc_data1[7]);
	soc_ethmac_crc32_checker_crc_next[2] <= (((((((((soc_ethmac_crc32_checker_crc_last[26] ^ soc_ethmac_crc32_checker_crc_data1[5]) ^ soc_ethmac_crc32_checker_crc_last[25]) ^ soc_ethmac_crc32_checker_crc_last[31]) ^ soc_ethmac_crc32_checker_crc_data1[0]) ^ soc_ethmac_crc32_checker_crc_data1[6]) ^ soc_ethmac_crc32_checker_crc_last[24]) ^ soc_ethmac_crc32_checker_crc_last[30]) ^ soc_ethmac_crc32_checker_crc_data1[1]) ^ soc_ethmac_crc32_checker_crc_data1[7]);
	soc_ethmac_crc32_checker_crc_next[3] <= (((((((soc_ethmac_crc32_checker_crc_last[27] ^ soc_ethmac_crc32_checker_crc_data1[4]) ^ soc_ethmac_crc32_checker_crc_last[26]) ^ soc_ethmac_crc32_checker_crc_data1[5]) ^ soc_ethmac_crc32_checker_crc_last[25]) ^ soc_ethmac_crc32_checker_crc_last[31]) ^ soc_ethmac_crc32_checker_crc_data1[0]) ^ soc_ethmac_crc32_checker_crc_data1[6]);
	soc_ethmac_crc32_checker_crc_next[4] <= (((((((((soc_ethmac_crc32_checker_crc_last[28] ^ soc_ethmac_crc32_checker_crc_data1[3]) ^ soc_ethmac_crc32_checker_crc_last[27]) ^ soc_ethmac_crc32_checker_crc_data1[4]) ^ soc_ethmac_crc32_checker_crc_last[26]) ^ soc_ethmac_crc32_checker_crc_data1[5]) ^ soc_ethmac_crc32_checker_crc_last[24]) ^ soc_ethmac_crc32_checker_crc_last[30]) ^ soc_ethmac_crc32_checker_crc_data1[1]) ^ soc_ethmac_crc32_checker_crc_data1[7]);
	soc_ethmac_crc32_checker_crc_next[5] <= (((((((((((((soc_ethmac_crc32_checker_crc_last[29] ^ soc_ethmac_crc32_checker_crc_data1[2]) ^ soc_ethmac_crc32_checker_crc_last[28]) ^ soc_ethmac_crc32_checker_crc_data1[3]) ^ soc_ethmac_crc32_checker_crc_last[27]) ^ soc_ethmac_crc32_checker_crc_data1[4]) ^ soc_ethmac_crc32_checker_crc_last[25]) ^ soc_ethmac_crc32_checker_crc_last[31]) ^ soc_ethmac_crc32_checker_crc_data1[0]) ^ soc_ethmac_crc32_checker_crc_data1[6]) ^ soc_ethmac_crc32_checker_crc_last[24]) ^ soc_ethmac_crc32_checker_crc_last[30]) ^ soc_ethmac_crc32_checker_crc_data1[1]) ^ soc_ethmac_crc32_checker_crc_data1[7]);
	soc_ethmac_crc32_checker_crc_next[6] <= (((((((((((soc_ethmac_crc32_checker_crc_last[30] ^ soc_ethmac_crc32_checker_crc_data1[1]) ^ soc_ethmac_crc32_checker_crc_last[29]) ^ soc_ethmac_crc32_checker_crc_data1[2]) ^ soc_ethmac_crc32_checker_crc_last[28]) ^ soc_ethmac_crc32_checker_crc_data1[3]) ^ soc_ethmac_crc32_checker_crc_last[26]) ^ soc_ethmac_crc32_checker_crc_data1[5]) ^ soc_ethmac_crc32_checker_crc_last[25]) ^ soc_ethmac_crc32_checker_crc_last[31]) ^ soc_ethmac_crc32_checker_crc_data1[0]) ^ soc_ethmac_crc32_checker_crc_data1[6]);
	soc_ethmac_crc32_checker_crc_next[7] <= (((((((((soc_ethmac_crc32_checker_crc_last[31] ^ soc_ethmac_crc32_checker_crc_data1[0]) ^ soc_ethmac_crc32_checker_crc_last[29]) ^ soc_ethmac_crc32_checker_crc_data1[2]) ^ soc_ethmac_crc32_checker_crc_last[27]) ^ soc_ethmac_crc32_checker_crc_data1[4]) ^ soc_ethmac_crc32_checker_crc_last[26]) ^ soc_ethmac_crc32_checker_crc_data1[5]) ^ soc_ethmac_crc32_checker_crc_last[24]) ^ soc_ethmac_crc32_checker_crc_data1[7]);
	soc_ethmac_crc32_checker_crc_next[8] <= ((((((((soc_ethmac_crc32_checker_crc_last[0] ^ soc_ethmac_crc32_checker_crc_last[28]) ^ soc_ethmac_crc32_checker_crc_data1[3]) ^ soc_ethmac_crc32_checker_crc_last[27]) ^ soc_ethmac_crc32_checker_crc_data1[4]) ^ soc_ethmac_crc32_checker_crc_last[25]) ^ soc_ethmac_crc32_checker_crc_data1[6]) ^ soc_ethmac_crc32_checker_crc_last[24]) ^ soc_ethmac_crc32_checker_crc_data1[7]);
	soc_ethmac_crc32_checker_crc_next[9] <= ((((((((soc_ethmac_crc32_checker_crc_last[1] ^ soc_ethmac_crc32_checker_crc_last[29]) ^ soc_ethmac_crc32_checker_crc_data1[2]) ^ soc_ethmac_crc32_checker_crc_last[28]) ^ soc_ethmac_crc32_checker_crc_data1[3]) ^ soc_ethmac_crc32_checker_crc_last[26]) ^ soc_ethmac_crc32_checker_crc_data1[5]) ^ soc_ethmac_crc32_checker_crc_last[25]) ^ soc_ethmac_crc32_checker_crc_data1[6]);
	soc_ethmac_crc32_checker_crc_next[10] <= ((((((((soc_ethmac_crc32_checker_crc_last[2] ^ soc_ethmac_crc32_checker_crc_last[29]) ^ soc_ethmac_crc32_checker_crc_data1[2]) ^ soc_ethmac_crc32_checker_crc_last[27]) ^ soc_ethmac_crc32_checker_crc_data1[4]) ^ soc_ethmac_crc32_checker_crc_last[26]) ^ soc_ethmac_crc32_checker_crc_data1[5]) ^ soc_ethmac_crc32_checker_crc_last[24]) ^ soc_ethmac_crc32_checker_crc_data1[7]);
	soc_ethmac_crc32_checker_crc_next[11] <= ((((((((soc_ethmac_crc32_checker_crc_last[3] ^ soc_ethmac_crc32_checker_crc_last[28]) ^ soc_ethmac_crc32_checker_crc_data1[3]) ^ soc_ethmac_crc32_checker_crc_last[27]) ^ soc_ethmac_crc32_checker_crc_data1[4]) ^ soc_ethmac_crc32_checker_crc_last[25]) ^ soc_ethmac_crc32_checker_crc_data1[6]) ^ soc_ethmac_crc32_checker_crc_last[24]) ^ soc_ethmac_crc32_checker_crc_data1[7]);
	soc_ethmac_crc32_checker_crc_next[12] <= ((((((((((((soc_ethmac_crc32_checker_crc_last[4] ^ soc_ethmac_crc32_checker_crc_last[29]) ^ soc_ethmac_crc32_checker_crc_data1[2]) ^ soc_ethmac_crc32_checker_crc_last[28]) ^ soc_ethmac_crc32_checker_crc_data1[3]) ^ soc_ethmac_crc32_checker_crc_last[26]) ^ soc_ethmac_crc32_checker_crc_data1[5]) ^ soc_ethmac_crc32_checker_crc_last[25]) ^ soc_ethmac_crc32_checker_crc_data1[6]) ^ soc_ethmac_crc32_checker_crc_last[24]) ^ soc_ethmac_crc32_checker_crc_last[30]) ^ soc_ethmac_crc32_checker_crc_data1[1]) ^ soc_ethmac_crc32_checker_crc_data1[7]);
	soc_ethmac_crc32_checker_crc_next[13] <= ((((((((((((soc_ethmac_crc32_checker_crc_last[5] ^ soc_ethmac_crc32_checker_crc_last[30]) ^ soc_ethmac_crc32_checker_crc_data1[1]) ^ soc_ethmac_crc32_checker_crc_last[29]) ^ soc_ethmac_crc32_checker_crc_data1[2]) ^ soc_ethmac_crc32_checker_crc_last[27]) ^ soc_ethmac_crc32_checker_crc_data1[4]) ^ soc_ethmac_crc32_checker_crc_last[26]) ^ soc_ethmac_crc32_checker_crc_data1[5]) ^ soc_ethmac_crc32_checker_crc_last[25]) ^ soc_ethmac_crc32_checker_crc_last[31]) ^ soc_ethmac_crc32_checker_crc_data1[0]) ^ soc_ethmac_crc32_checker_crc_data1[6]);
	soc_ethmac_crc32_checker_crc_next[14] <= ((((((((((soc_ethmac_crc32_checker_crc_last[6] ^ soc_ethmac_crc32_checker_crc_last[31]) ^ soc_ethmac_crc32_checker_crc_data1[0]) ^ soc_ethmac_crc32_checker_crc_last[30]) ^ soc_ethmac_crc32_checker_crc_data1[1]) ^ soc_ethmac_crc32_checker_crc_last[28]) ^ soc_ethmac_crc32_checker_crc_data1[3]) ^ soc_ethmac_crc32_checker_crc_last[27]) ^ soc_ethmac_crc32_checker_crc_data1[4]) ^ soc_ethmac_crc32_checker_crc_last[26]) ^ soc_ethmac_crc32_checker_crc_data1[5]);
	soc_ethmac_crc32_checker_crc_next[15] <= ((((((((soc_ethmac_crc32_checker_crc_last[7] ^ soc_ethmac_crc32_checker_crc_last[31]) ^ soc_ethmac_crc32_checker_crc_data1[0]) ^ soc_ethmac_crc32_checker_crc_last[29]) ^ soc_ethmac_crc32_checker_crc_data1[2]) ^ soc_ethmac_crc32_checker_crc_last[28]) ^ soc_ethmac_crc32_checker_crc_data1[3]) ^ soc_ethmac_crc32_checker_crc_last[27]) ^ soc_ethmac_crc32_checker_crc_data1[4]);
	soc_ethmac_crc32_checker_crc_next[16] <= ((((((soc_ethmac_crc32_checker_crc_last[8] ^ soc_ethmac_crc32_checker_crc_last[29]) ^ soc_ethmac_crc32_checker_crc_data1[2]) ^ soc_ethmac_crc32_checker_crc_last[28]) ^ soc_ethmac_crc32_checker_crc_data1[3]) ^ soc_ethmac_crc32_checker_crc_last[24]) ^ soc_ethmac_crc32_checker_crc_data1[7]);
	soc_ethmac_crc32_checker_crc_next[17] <= ((((((soc_ethmac_crc32_checker_crc_last[9] ^ soc_ethmac_crc32_checker_crc_last[30]) ^ soc_ethmac_crc32_checker_crc_data1[1]) ^ soc_ethmac_crc32_checker_crc_last[29]) ^ soc_ethmac_crc32_checker_crc_data1[2]) ^ soc_ethmac_crc32_checker_crc_last[25]) ^ soc_ethmac_crc32_checker_crc_data1[6]);
	soc_ethmac_crc32_checker_crc_next[18] <= ((((((soc_ethmac_crc32_checker_crc_last[10] ^ soc_ethmac_crc32_checker_crc_last[31]) ^ soc_ethmac_crc32_checker_crc_data1[0]) ^ soc_ethmac_crc32_checker_crc_last[30]) ^ soc_ethmac_crc32_checker_crc_data1[1]) ^ soc_ethmac_crc32_checker_crc_last[26]) ^ soc_ethmac_crc32_checker_crc_data1[5]);
	soc_ethmac_crc32_checker_crc_next[19] <= ((((soc_ethmac_crc32_checker_crc_last[11] ^ soc_ethmac_crc32_checker_crc_last[31]) ^ soc_ethmac_crc32_checker_crc_data1[0]) ^ soc_ethmac_crc32_checker_crc_last[27]) ^ soc_ethmac_crc32_checker_crc_data1[4]);
	soc_ethmac_crc32_checker_crc_next[20] <= ((soc_ethmac_crc32_checker_crc_last[12] ^ soc_ethmac_crc32_checker_crc_last[28]) ^ soc_ethmac_crc32_checker_crc_data1[3]);
	soc_ethmac_crc32_checker_crc_next[21] <= ((soc_ethmac_crc32_checker_crc_last[13] ^ soc_ethmac_crc32_checker_crc_last[29]) ^ soc_ethmac_crc32_checker_crc_data1[2]);
	soc_ethmac_crc32_checker_crc_next[22] <= ((soc_ethmac_crc32_checker_crc_last[14] ^ soc_ethmac_crc32_checker_crc_last[24]) ^ soc_ethmac_crc32_checker_crc_data1[7]);
	soc_ethmac_crc32_checker_crc_next[23] <= ((((((soc_ethmac_crc32_checker_crc_last[15] ^ soc_ethmac_crc32_checker_crc_last[25]) ^ soc_ethmac_crc32_checker_crc_data1[6]) ^ soc_ethmac_crc32_checker_crc_last[24]) ^ soc_ethmac_crc32_checker_crc_last[30]) ^ soc_ethmac_crc32_checker_crc_data1[1]) ^ soc_ethmac_crc32_checker_crc_data1[7]);
	soc_ethmac_crc32_checker_crc_next[24] <= ((((((soc_ethmac_crc32_checker_crc_last[16] ^ soc_ethmac_crc32_checker_crc_last[26]) ^ soc_ethmac_crc32_checker_crc_data1[5]) ^ soc_ethmac_crc32_checker_crc_last[25]) ^ soc_ethmac_crc32_checker_crc_last[31]) ^ soc_ethmac_crc32_checker_crc_data1[0]) ^ soc_ethmac_crc32_checker_crc_data1[6]);
	soc_ethmac_crc32_checker_crc_next[25] <= ((((soc_ethmac_crc32_checker_crc_last[17] ^ soc_ethmac_crc32_checker_crc_last[27]) ^ soc_ethmac_crc32_checker_crc_data1[4]) ^ soc_ethmac_crc32_checker_crc_last[26]) ^ soc_ethmac_crc32_checker_crc_data1[5]);
	soc_ethmac_crc32_checker_crc_next[26] <= ((((((((soc_ethmac_crc32_checker_crc_last[18] ^ soc_ethmac_crc32_checker_crc_last[28]) ^ soc_ethmac_crc32_checker_crc_data1[3]) ^ soc_ethmac_crc32_checker_crc_last[27]) ^ soc_ethmac_crc32_checker_crc_data1[4]) ^ soc_ethmac_crc32_checker_crc_last[24]) ^ soc_ethmac_crc32_checker_crc_last[30]) ^ soc_ethmac_crc32_checker_crc_data1[1]) ^ soc_ethmac_crc32_checker_crc_data1[7]);
	soc_ethmac_crc32_checker_crc_next[27] <= ((((((((soc_ethmac_crc32_checker_crc_last[19] ^ soc_ethmac_crc32_checker_crc_last[29]) ^ soc_ethmac_crc32_checker_crc_data1[2]) ^ soc_ethmac_crc32_checker_crc_last[28]) ^ soc_ethmac_crc32_checker_crc_data1[3]) ^ soc_ethmac_crc32_checker_crc_last[25]) ^ soc_ethmac_crc32_checker_crc_last[31]) ^ soc_ethmac_crc32_checker_crc_data1[0]) ^ soc_ethmac_crc32_checker_crc_data1[6]);
	soc_ethmac_crc32_checker_crc_next[28] <= ((((((soc_ethmac_crc32_checker_crc_last[20] ^ soc_ethmac_crc32_checker_crc_last[30]) ^ soc_ethmac_crc32_checker_crc_data1[1]) ^ soc_ethmac_crc32_checker_crc_last[29]) ^ soc_ethmac_crc32_checker_crc_data1[2]) ^ soc_ethmac_crc32_checker_crc_last[26]) ^ soc_ethmac_crc32_checker_crc_data1[5]);
	soc_ethmac_crc32_checker_crc_next[29] <= ((((((soc_ethmac_crc32_checker_crc_last[21] ^ soc_ethmac_crc32_checker_crc_last[31]) ^ soc_ethmac_crc32_checker_crc_data1[0]) ^ soc_ethmac_crc32_checker_crc_last[30]) ^ soc_ethmac_crc32_checker_crc_data1[1]) ^ soc_ethmac_crc32_checker_crc_last[27]) ^ soc_ethmac_crc32_checker_crc_data1[4]);
	soc_ethmac_crc32_checker_crc_next[30] <= ((((soc_ethmac_crc32_checker_crc_last[22] ^ soc_ethmac_crc32_checker_crc_last[31]) ^ soc_ethmac_crc32_checker_crc_data1[0]) ^ soc_ethmac_crc32_checker_crc_last[28]) ^ soc_ethmac_crc32_checker_crc_data1[3]);
	soc_ethmac_crc32_checker_crc_next[31] <= ((soc_ethmac_crc32_checker_crc_last[23] ^ soc_ethmac_crc32_checker_crc_last[29]) ^ soc_ethmac_crc32_checker_crc_data1[2]);
end
assign soc_ethmac_crc32_checker_syncfifo_syncfifo_din = {soc_ethmac_crc32_checker_syncfifo_fifo_in_last, soc_ethmac_crc32_checker_syncfifo_fifo_in_first, soc_ethmac_crc32_checker_syncfifo_fifo_in_payload_error, soc_ethmac_crc32_checker_syncfifo_fifo_in_payload_last_be, soc_ethmac_crc32_checker_syncfifo_fifo_in_payload_data};
assign {soc_ethmac_crc32_checker_syncfifo_fifo_out_last, soc_ethmac_crc32_checker_syncfifo_fifo_out_first, soc_ethmac_crc32_checker_syncfifo_fifo_out_payload_error, soc_ethmac_crc32_checker_syncfifo_fifo_out_payload_last_be, soc_ethmac_crc32_checker_syncfifo_fifo_out_payload_data} = soc_ethmac_crc32_checker_syncfifo_syncfifo_dout;
assign soc_ethmac_crc32_checker_syncfifo_sink_ready = soc_ethmac_crc32_checker_syncfifo_syncfifo_writable;
assign soc_ethmac_crc32_checker_syncfifo_syncfifo_we = soc_ethmac_crc32_checker_syncfifo_sink_valid;
assign soc_ethmac_crc32_checker_syncfifo_fifo_in_first = soc_ethmac_crc32_checker_syncfifo_sink_first;
assign soc_ethmac_crc32_checker_syncfifo_fifo_in_last = soc_ethmac_crc32_checker_syncfifo_sink_last;
assign soc_ethmac_crc32_checker_syncfifo_fifo_in_payload_data = soc_ethmac_crc32_checker_syncfifo_sink_payload_data;
assign soc_ethmac_crc32_checker_syncfifo_fifo_in_payload_last_be = soc_ethmac_crc32_checker_syncfifo_sink_payload_last_be;
assign soc_ethmac_crc32_checker_syncfifo_fifo_in_payload_error = soc_ethmac_crc32_checker_syncfifo_sink_payload_error;
assign soc_ethmac_crc32_checker_syncfifo_source_valid = soc_ethmac_crc32_checker_syncfifo_syncfifo_readable;
assign soc_ethmac_crc32_checker_syncfifo_source_first = soc_ethmac_crc32_checker_syncfifo_fifo_out_first;
assign soc_ethmac_crc32_checker_syncfifo_source_last = soc_ethmac_crc32_checker_syncfifo_fifo_out_last;
assign soc_ethmac_crc32_checker_syncfifo_source_payload_data = soc_ethmac_crc32_checker_syncfifo_fifo_out_payload_data;
assign soc_ethmac_crc32_checker_syncfifo_source_payload_last_be = soc_ethmac_crc32_checker_syncfifo_fifo_out_payload_last_be;
assign soc_ethmac_crc32_checker_syncfifo_source_payload_error = soc_ethmac_crc32_checker_syncfifo_fifo_out_payload_error;
assign soc_ethmac_crc32_checker_syncfifo_syncfifo_re = soc_ethmac_crc32_checker_syncfifo_source_ready;
always @(*) begin
	soc_ethmac_crc32_checker_syncfifo_wrport_adr <= 3'd0;
	if (soc_ethmac_crc32_checker_syncfifo_replace) begin
		soc_ethmac_crc32_checker_syncfifo_wrport_adr <= (soc_ethmac_crc32_checker_syncfifo_produce - 1'd1);
	end else begin
		soc_ethmac_crc32_checker_syncfifo_wrport_adr <= soc_ethmac_crc32_checker_syncfifo_produce;
	end
end
assign soc_ethmac_crc32_checker_syncfifo_wrport_dat_w = soc_ethmac_crc32_checker_syncfifo_syncfifo_din;
assign soc_ethmac_crc32_checker_syncfifo_wrport_we = (soc_ethmac_crc32_checker_syncfifo_syncfifo_we & (soc_ethmac_crc32_checker_syncfifo_syncfifo_writable | soc_ethmac_crc32_checker_syncfifo_replace));
assign soc_ethmac_crc32_checker_syncfifo_do_read = (soc_ethmac_crc32_checker_syncfifo_syncfifo_readable & soc_ethmac_crc32_checker_syncfifo_syncfifo_re);
assign soc_ethmac_crc32_checker_syncfifo_rdport_adr = soc_ethmac_crc32_checker_syncfifo_consume;
assign soc_ethmac_crc32_checker_syncfifo_syncfifo_dout = soc_ethmac_crc32_checker_syncfifo_rdport_dat_r;
assign soc_ethmac_crc32_checker_syncfifo_syncfifo_writable = (soc_ethmac_crc32_checker_syncfifo_level != 3'd5);
assign soc_ethmac_crc32_checker_syncfifo_syncfifo_readable = (soc_ethmac_crc32_checker_syncfifo_level != 1'd0);
always @(*) begin
	soc_ethmac_crc32_checker_crc_ce <= 1'd0;
	soc_ethmac_crc32_checker_fifo_reset <= 1'd0;
	vns_clockdomainsrenamer5_next_state <= 2'd0;
	soc_ethmac_crc32_checker_crc_reset <= 1'd0;
	vns_clockdomainsrenamer5_next_state <= vns_clockdomainsrenamer5_state;
	case (vns_clockdomainsrenamer5_state)
		1'd1: begin
			if ((soc_ethmac_crc32_checker_sink_sink_valid & soc_ethmac_crc32_checker_sink_sink_ready)) begin
				soc_ethmac_crc32_checker_crc_ce <= 1'd1;
				vns_clockdomainsrenamer5_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if ((soc_ethmac_crc32_checker_sink_sink_valid & soc_ethmac_crc32_checker_sink_sink_ready)) begin
				soc_ethmac_crc32_checker_crc_ce <= 1'd1;
				if (soc_ethmac_crc32_checker_sink_sink_last) begin
					vns_clockdomainsrenamer5_next_state <= 1'd0;
				end
			end
		end
		default: begin
			soc_ethmac_crc32_checker_crc_reset <= 1'd1;
			soc_ethmac_crc32_checker_fifo_reset <= 1'd1;
			vns_clockdomainsrenamer5_next_state <= 1'd1;
		end
	endcase
end
assign soc_ethmac_padding_inserter_counter_done = (soc_ethmac_padding_inserter_counter >= 6'd59);
always @(*) begin
	soc_ethmac_padding_inserter_source_valid <= 1'd0;
	vns_clockdomainsrenamer6_next_state <= 1'd0;
	soc_ethmac_padding_inserter_source_first <= 1'd0;
	soc_ethmac_padding_inserter_source_last <= 1'd0;
	soc_ethmac_padding_inserter_source_payload_data <= 8'd0;
	soc_ethmac_padding_inserter_source_payload_last_be <= 1'd0;
	soc_ethmac_padding_inserter_source_payload_error <= 1'd0;
	soc_ethmac_padding_inserter_counter_reset <= 1'd0;
	soc_ethmac_padding_inserter_counter_ce <= 1'd0;
	soc_ethmac_padding_inserter_sink_ready <= 1'd0;
	vns_clockdomainsrenamer6_next_state <= vns_clockdomainsrenamer6_state;
	case (vns_clockdomainsrenamer6_state)
		1'd1: begin
			soc_ethmac_padding_inserter_source_valid <= 1'd1;
			soc_ethmac_padding_inserter_source_last <= soc_ethmac_padding_inserter_counter_done;
			soc_ethmac_padding_inserter_source_payload_data <= 1'd0;
			if ((soc_ethmac_padding_inserter_source_valid & soc_ethmac_padding_inserter_source_ready)) begin
				soc_ethmac_padding_inserter_counter_ce <= 1'd1;
				if (soc_ethmac_padding_inserter_counter_done) begin
					soc_ethmac_padding_inserter_counter_reset <= 1'd1;
					vns_clockdomainsrenamer6_next_state <= 1'd0;
				end
			end
		end
		default: begin
			soc_ethmac_padding_inserter_source_valid <= soc_ethmac_padding_inserter_sink_valid;
			soc_ethmac_padding_inserter_sink_ready <= soc_ethmac_padding_inserter_source_ready;
			soc_ethmac_padding_inserter_source_first <= soc_ethmac_padding_inserter_sink_first;
			soc_ethmac_padding_inserter_source_last <= soc_ethmac_padding_inserter_sink_last;
			soc_ethmac_padding_inserter_source_payload_data <= soc_ethmac_padding_inserter_sink_payload_data;
			soc_ethmac_padding_inserter_source_payload_last_be <= soc_ethmac_padding_inserter_sink_payload_last_be;
			soc_ethmac_padding_inserter_source_payload_error <= soc_ethmac_padding_inserter_sink_payload_error;
			if ((soc_ethmac_padding_inserter_source_valid & soc_ethmac_padding_inserter_source_ready)) begin
				soc_ethmac_padding_inserter_counter_ce <= 1'd1;
				if (soc_ethmac_padding_inserter_sink_last) begin
					if ((~soc_ethmac_padding_inserter_counter_done)) begin
						soc_ethmac_padding_inserter_source_last <= 1'd0;
						vns_clockdomainsrenamer6_next_state <= 1'd1;
					end else begin
						soc_ethmac_padding_inserter_counter_reset <= 1'd1;
					end
				end
			end
		end
	endcase
end
assign soc_ethmac_padding_checker_source_valid = soc_ethmac_padding_checker_sink_valid;
assign soc_ethmac_padding_checker_sink_ready = soc_ethmac_padding_checker_source_ready;
assign soc_ethmac_padding_checker_source_first = soc_ethmac_padding_checker_sink_first;
assign soc_ethmac_padding_checker_source_last = soc_ethmac_padding_checker_sink_last;
assign soc_ethmac_padding_checker_source_payload_data = soc_ethmac_padding_checker_sink_payload_data;
assign soc_ethmac_padding_checker_source_payload_last_be = soc_ethmac_padding_checker_sink_payload_last_be;
assign soc_ethmac_padding_checker_source_payload_error = soc_ethmac_padding_checker_sink_payload_error;
assign soc_ethmac_tx_last_be_source_valid = (soc_ethmac_tx_last_be_sink_valid & soc_ethmac_tx_last_be_ongoing);
assign soc_ethmac_tx_last_be_source_last = soc_ethmac_tx_last_be_sink_payload_last_be;
assign soc_ethmac_tx_last_be_source_payload_data = soc_ethmac_tx_last_be_sink_payload_data;
assign soc_ethmac_tx_last_be_sink_ready = soc_ethmac_tx_last_be_source_ready;
assign soc_ethmac_rx_last_be_source_valid = soc_ethmac_rx_last_be_sink_valid;
assign soc_ethmac_rx_last_be_sink_ready = soc_ethmac_rx_last_be_source_ready;
assign soc_ethmac_rx_last_be_source_first = soc_ethmac_rx_last_be_sink_first;
assign soc_ethmac_rx_last_be_source_last = soc_ethmac_rx_last_be_sink_last;
assign soc_ethmac_rx_last_be_source_payload_data = soc_ethmac_rx_last_be_sink_payload_data;
assign soc_ethmac_rx_last_be_source_payload_error = soc_ethmac_rx_last_be_sink_payload_error;
always @(*) begin
	soc_ethmac_rx_last_be_source_payload_last_be <= 1'd0;
	soc_ethmac_rx_last_be_source_payload_last_be <= soc_ethmac_rx_last_be_sink_payload_last_be;
	soc_ethmac_rx_last_be_source_payload_last_be <= soc_ethmac_rx_last_be_sink_last;
end
assign soc_ethmac_tx_converter_converter_sink_valid = soc_ethmac_tx_converter_sink_valid;
assign soc_ethmac_tx_converter_converter_sink_first = soc_ethmac_tx_converter_sink_first;
assign soc_ethmac_tx_converter_converter_sink_last = soc_ethmac_tx_converter_sink_last;
assign soc_ethmac_tx_converter_sink_ready = soc_ethmac_tx_converter_converter_sink_ready;
always @(*) begin
	soc_ethmac_tx_converter_converter_sink_payload_data <= 40'd0;
	soc_ethmac_tx_converter_converter_sink_payload_data[7:0] <= soc_ethmac_tx_converter_sink_payload_data[7:0];
	soc_ethmac_tx_converter_converter_sink_payload_data[8] <= soc_ethmac_tx_converter_sink_payload_last_be[0];
	soc_ethmac_tx_converter_converter_sink_payload_data[9] <= soc_ethmac_tx_converter_sink_payload_error[0];
	soc_ethmac_tx_converter_converter_sink_payload_data[17:10] <= soc_ethmac_tx_converter_sink_payload_data[15:8];
	soc_ethmac_tx_converter_converter_sink_payload_data[18] <= soc_ethmac_tx_converter_sink_payload_last_be[1];
	soc_ethmac_tx_converter_converter_sink_payload_data[19] <= soc_ethmac_tx_converter_sink_payload_error[1];
	soc_ethmac_tx_converter_converter_sink_payload_data[27:20] <= soc_ethmac_tx_converter_sink_payload_data[23:16];
	soc_ethmac_tx_converter_converter_sink_payload_data[28] <= soc_ethmac_tx_converter_sink_payload_last_be[2];
	soc_ethmac_tx_converter_converter_sink_payload_data[29] <= soc_ethmac_tx_converter_sink_payload_error[2];
	soc_ethmac_tx_converter_converter_sink_payload_data[37:30] <= soc_ethmac_tx_converter_sink_payload_data[31:24];
	soc_ethmac_tx_converter_converter_sink_payload_data[38] <= soc_ethmac_tx_converter_sink_payload_last_be[3];
	soc_ethmac_tx_converter_converter_sink_payload_data[39] <= soc_ethmac_tx_converter_sink_payload_error[3];
end
assign soc_ethmac_tx_converter_source_valid = soc_ethmac_tx_converter_source_source_valid;
assign soc_ethmac_tx_converter_source_first = soc_ethmac_tx_converter_source_source_first;
assign soc_ethmac_tx_converter_source_last = soc_ethmac_tx_converter_source_source_last;
assign soc_ethmac_tx_converter_source_source_ready = soc_ethmac_tx_converter_source_ready;
assign {soc_ethmac_tx_converter_source_payload_error, soc_ethmac_tx_converter_source_payload_last_be, soc_ethmac_tx_converter_source_payload_data} = soc_ethmac_tx_converter_source_source_payload_data;
assign soc_ethmac_tx_converter_source_source_valid = soc_ethmac_tx_converter_converter_source_valid;
assign soc_ethmac_tx_converter_converter_source_ready = soc_ethmac_tx_converter_source_source_ready;
assign soc_ethmac_tx_converter_source_source_first = soc_ethmac_tx_converter_converter_source_first;
assign soc_ethmac_tx_converter_source_source_last = soc_ethmac_tx_converter_converter_source_last;
assign soc_ethmac_tx_converter_source_source_payload_data = soc_ethmac_tx_converter_converter_source_payload_data;
assign soc_ethmac_tx_converter_converter_first = (soc_ethmac_tx_converter_converter_mux == 1'd0);
assign soc_ethmac_tx_converter_converter_last = (soc_ethmac_tx_converter_converter_mux == 2'd3);
assign soc_ethmac_tx_converter_converter_source_valid = soc_ethmac_tx_converter_converter_sink_valid;
assign soc_ethmac_tx_converter_converter_source_first = (soc_ethmac_tx_converter_converter_sink_first & soc_ethmac_tx_converter_converter_first);
assign soc_ethmac_tx_converter_converter_source_last = (soc_ethmac_tx_converter_converter_sink_last & soc_ethmac_tx_converter_converter_last);
assign soc_ethmac_tx_converter_converter_sink_ready = (soc_ethmac_tx_converter_converter_last & soc_ethmac_tx_converter_converter_source_ready);
always @(*) begin
	soc_ethmac_tx_converter_converter_source_payload_data <= 10'd0;
	case (soc_ethmac_tx_converter_converter_mux)
		1'd0: begin
			soc_ethmac_tx_converter_converter_source_payload_data <= soc_ethmac_tx_converter_converter_sink_payload_data[39:30];
		end
		1'd1: begin
			soc_ethmac_tx_converter_converter_source_payload_data <= soc_ethmac_tx_converter_converter_sink_payload_data[29:20];
		end
		2'd2: begin
			soc_ethmac_tx_converter_converter_source_payload_data <= soc_ethmac_tx_converter_converter_sink_payload_data[19:10];
		end
		default: begin
			soc_ethmac_tx_converter_converter_source_payload_data <= soc_ethmac_tx_converter_converter_sink_payload_data[9:0];
		end
	endcase
end
assign soc_ethmac_tx_converter_converter_source_payload_valid_token_count = soc_ethmac_tx_converter_converter_last;
assign soc_ethmac_rx_converter_converter_sink_valid = soc_ethmac_rx_converter_sink_valid;
assign soc_ethmac_rx_converter_converter_sink_first = soc_ethmac_rx_converter_sink_first;
assign soc_ethmac_rx_converter_converter_sink_last = soc_ethmac_rx_converter_sink_last;
assign soc_ethmac_rx_converter_sink_ready = soc_ethmac_rx_converter_converter_sink_ready;
assign soc_ethmac_rx_converter_converter_sink_payload_data = {soc_ethmac_rx_converter_sink_payload_error, soc_ethmac_rx_converter_sink_payload_last_be, soc_ethmac_rx_converter_sink_payload_data};
assign soc_ethmac_rx_converter_source_valid = soc_ethmac_rx_converter_source_source_valid;
assign soc_ethmac_rx_converter_source_first = soc_ethmac_rx_converter_source_source_first;
assign soc_ethmac_rx_converter_source_last = soc_ethmac_rx_converter_source_source_last;
assign soc_ethmac_rx_converter_source_source_ready = soc_ethmac_rx_converter_source_ready;
always @(*) begin
	soc_ethmac_rx_converter_source_payload_data <= 32'd0;
	soc_ethmac_rx_converter_source_payload_data[7:0] <= soc_ethmac_rx_converter_source_source_payload_data[7:0];
	soc_ethmac_rx_converter_source_payload_data[15:8] <= soc_ethmac_rx_converter_source_source_payload_data[17:10];
	soc_ethmac_rx_converter_source_payload_data[23:16] <= soc_ethmac_rx_converter_source_source_payload_data[27:20];
	soc_ethmac_rx_converter_source_payload_data[31:24] <= soc_ethmac_rx_converter_source_source_payload_data[37:30];
end
always @(*) begin
	soc_ethmac_rx_converter_source_payload_last_be <= 4'd0;
	soc_ethmac_rx_converter_source_payload_last_be[0] <= soc_ethmac_rx_converter_source_source_payload_data[8];
	soc_ethmac_rx_converter_source_payload_last_be[1] <= soc_ethmac_rx_converter_source_source_payload_data[18];
	soc_ethmac_rx_converter_source_payload_last_be[2] <= soc_ethmac_rx_converter_source_source_payload_data[28];
	soc_ethmac_rx_converter_source_payload_last_be[3] <= soc_ethmac_rx_converter_source_source_payload_data[38];
end
always @(*) begin
	soc_ethmac_rx_converter_source_payload_error <= 4'd0;
	soc_ethmac_rx_converter_source_payload_error[0] <= soc_ethmac_rx_converter_source_source_payload_data[9];
	soc_ethmac_rx_converter_source_payload_error[1] <= soc_ethmac_rx_converter_source_source_payload_data[19];
	soc_ethmac_rx_converter_source_payload_error[2] <= soc_ethmac_rx_converter_source_source_payload_data[29];
	soc_ethmac_rx_converter_source_payload_error[3] <= soc_ethmac_rx_converter_source_source_payload_data[39];
end
assign soc_ethmac_rx_converter_source_source_valid = soc_ethmac_rx_converter_converter_source_valid;
assign soc_ethmac_rx_converter_converter_source_ready = soc_ethmac_rx_converter_source_source_ready;
assign soc_ethmac_rx_converter_source_source_first = soc_ethmac_rx_converter_converter_source_first;
assign soc_ethmac_rx_converter_source_source_last = soc_ethmac_rx_converter_converter_source_last;
assign soc_ethmac_rx_converter_source_source_payload_data = soc_ethmac_rx_converter_converter_source_payload_data;
assign soc_ethmac_rx_converter_converter_sink_ready = ((~soc_ethmac_rx_converter_converter_strobe_all) | soc_ethmac_rx_converter_converter_source_ready);
assign soc_ethmac_rx_converter_converter_source_valid = soc_ethmac_rx_converter_converter_strobe_all;
assign soc_ethmac_rx_converter_converter_load_part = (soc_ethmac_rx_converter_converter_sink_valid & soc_ethmac_rx_converter_converter_sink_ready);
assign soc_ethmac_tx_cdc_asyncfifo_din = {soc_ethmac_tx_cdc_fifo_in_last, soc_ethmac_tx_cdc_fifo_in_first, soc_ethmac_tx_cdc_fifo_in_payload_error, soc_ethmac_tx_cdc_fifo_in_payload_last_be, soc_ethmac_tx_cdc_fifo_in_payload_data};
assign {soc_ethmac_tx_cdc_fifo_out_last, soc_ethmac_tx_cdc_fifo_out_first, soc_ethmac_tx_cdc_fifo_out_payload_error, soc_ethmac_tx_cdc_fifo_out_payload_last_be, soc_ethmac_tx_cdc_fifo_out_payload_data} = soc_ethmac_tx_cdc_asyncfifo_dout;
assign soc_ethmac_tx_cdc_sink_ready = soc_ethmac_tx_cdc_asyncfifo_writable;
assign soc_ethmac_tx_cdc_asyncfifo_we = soc_ethmac_tx_cdc_sink_valid;
assign soc_ethmac_tx_cdc_fifo_in_first = soc_ethmac_tx_cdc_sink_first;
assign soc_ethmac_tx_cdc_fifo_in_last = soc_ethmac_tx_cdc_sink_last;
assign soc_ethmac_tx_cdc_fifo_in_payload_data = soc_ethmac_tx_cdc_sink_payload_data;
assign soc_ethmac_tx_cdc_fifo_in_payload_last_be = soc_ethmac_tx_cdc_sink_payload_last_be;
assign soc_ethmac_tx_cdc_fifo_in_payload_error = soc_ethmac_tx_cdc_sink_payload_error;
assign soc_ethmac_tx_cdc_source_valid = soc_ethmac_tx_cdc_asyncfifo_readable;
assign soc_ethmac_tx_cdc_source_first = soc_ethmac_tx_cdc_fifo_out_first;
assign soc_ethmac_tx_cdc_source_last = soc_ethmac_tx_cdc_fifo_out_last;
assign soc_ethmac_tx_cdc_source_payload_data = soc_ethmac_tx_cdc_fifo_out_payload_data;
assign soc_ethmac_tx_cdc_source_payload_last_be = soc_ethmac_tx_cdc_fifo_out_payload_last_be;
assign soc_ethmac_tx_cdc_source_payload_error = soc_ethmac_tx_cdc_fifo_out_payload_error;
assign soc_ethmac_tx_cdc_asyncfifo_re = soc_ethmac_tx_cdc_source_ready;
assign soc_ethmac_tx_cdc_graycounter0_ce = (soc_ethmac_tx_cdc_asyncfifo_writable & soc_ethmac_tx_cdc_asyncfifo_we);
assign soc_ethmac_tx_cdc_graycounter1_ce = (soc_ethmac_tx_cdc_asyncfifo_readable & soc_ethmac_tx_cdc_asyncfifo_re);
assign soc_ethmac_tx_cdc_asyncfifo_writable = (((soc_ethmac_tx_cdc_graycounter0_q[6] == soc_ethmac_tx_cdc_consume_wdomain[6]) | (soc_ethmac_tx_cdc_graycounter0_q[5] == soc_ethmac_tx_cdc_consume_wdomain[5])) | (soc_ethmac_tx_cdc_graycounter0_q[4:0] != soc_ethmac_tx_cdc_consume_wdomain[4:0]));
assign soc_ethmac_tx_cdc_asyncfifo_readable = (soc_ethmac_tx_cdc_graycounter1_q != soc_ethmac_tx_cdc_produce_rdomain);
assign soc_ethmac_tx_cdc_wrport_adr = soc_ethmac_tx_cdc_graycounter0_q_binary[5:0];
assign soc_ethmac_tx_cdc_wrport_dat_w = soc_ethmac_tx_cdc_asyncfifo_din;
assign soc_ethmac_tx_cdc_wrport_we = soc_ethmac_tx_cdc_graycounter0_ce;
assign soc_ethmac_tx_cdc_rdport_adr = soc_ethmac_tx_cdc_graycounter1_q_next_binary[5:0];
assign soc_ethmac_tx_cdc_asyncfifo_dout = soc_ethmac_tx_cdc_rdport_dat_r;
always @(*) begin
	soc_ethmac_tx_cdc_graycounter0_q_next_binary <= 7'd0;
	if (soc_ethmac_tx_cdc_graycounter0_ce) begin
		soc_ethmac_tx_cdc_graycounter0_q_next_binary <= (soc_ethmac_tx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		soc_ethmac_tx_cdc_graycounter0_q_next_binary <= soc_ethmac_tx_cdc_graycounter0_q_binary;
	end
end
assign soc_ethmac_tx_cdc_graycounter0_q_next = (soc_ethmac_tx_cdc_graycounter0_q_next_binary ^ soc_ethmac_tx_cdc_graycounter0_q_next_binary[6:1]);
always @(*) begin
	soc_ethmac_tx_cdc_graycounter1_q_next_binary <= 7'd0;
	if (soc_ethmac_tx_cdc_graycounter1_ce) begin
		soc_ethmac_tx_cdc_graycounter1_q_next_binary <= (soc_ethmac_tx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		soc_ethmac_tx_cdc_graycounter1_q_next_binary <= soc_ethmac_tx_cdc_graycounter1_q_binary;
	end
end
assign soc_ethmac_tx_cdc_graycounter1_q_next = (soc_ethmac_tx_cdc_graycounter1_q_next_binary ^ soc_ethmac_tx_cdc_graycounter1_q_next_binary[6:1]);
assign soc_ethmac_rx_cdc_asyncfifo_din = {soc_ethmac_rx_cdc_fifo_in_last, soc_ethmac_rx_cdc_fifo_in_first, soc_ethmac_rx_cdc_fifo_in_payload_error, soc_ethmac_rx_cdc_fifo_in_payload_last_be, soc_ethmac_rx_cdc_fifo_in_payload_data};
assign {soc_ethmac_rx_cdc_fifo_out_last, soc_ethmac_rx_cdc_fifo_out_first, soc_ethmac_rx_cdc_fifo_out_payload_error, soc_ethmac_rx_cdc_fifo_out_payload_last_be, soc_ethmac_rx_cdc_fifo_out_payload_data} = soc_ethmac_rx_cdc_asyncfifo_dout;
assign soc_ethmac_rx_cdc_sink_ready = soc_ethmac_rx_cdc_asyncfifo_writable;
assign soc_ethmac_rx_cdc_asyncfifo_we = soc_ethmac_rx_cdc_sink_valid;
assign soc_ethmac_rx_cdc_fifo_in_first = soc_ethmac_rx_cdc_sink_first;
assign soc_ethmac_rx_cdc_fifo_in_last = soc_ethmac_rx_cdc_sink_last;
assign soc_ethmac_rx_cdc_fifo_in_payload_data = soc_ethmac_rx_cdc_sink_payload_data;
assign soc_ethmac_rx_cdc_fifo_in_payload_last_be = soc_ethmac_rx_cdc_sink_payload_last_be;
assign soc_ethmac_rx_cdc_fifo_in_payload_error = soc_ethmac_rx_cdc_sink_payload_error;
assign soc_ethmac_rx_cdc_source_valid = soc_ethmac_rx_cdc_asyncfifo_readable;
assign soc_ethmac_rx_cdc_source_first = soc_ethmac_rx_cdc_fifo_out_first;
assign soc_ethmac_rx_cdc_source_last = soc_ethmac_rx_cdc_fifo_out_last;
assign soc_ethmac_rx_cdc_source_payload_data = soc_ethmac_rx_cdc_fifo_out_payload_data;
assign soc_ethmac_rx_cdc_source_payload_last_be = soc_ethmac_rx_cdc_fifo_out_payload_last_be;
assign soc_ethmac_rx_cdc_source_payload_error = soc_ethmac_rx_cdc_fifo_out_payload_error;
assign soc_ethmac_rx_cdc_asyncfifo_re = soc_ethmac_rx_cdc_source_ready;
assign soc_ethmac_rx_cdc_graycounter0_ce = (soc_ethmac_rx_cdc_asyncfifo_writable & soc_ethmac_rx_cdc_asyncfifo_we);
assign soc_ethmac_rx_cdc_graycounter1_ce = (soc_ethmac_rx_cdc_asyncfifo_readable & soc_ethmac_rx_cdc_asyncfifo_re);
assign soc_ethmac_rx_cdc_asyncfifo_writable = (((soc_ethmac_rx_cdc_graycounter0_q[6] == soc_ethmac_rx_cdc_consume_wdomain[6]) | (soc_ethmac_rx_cdc_graycounter0_q[5] == soc_ethmac_rx_cdc_consume_wdomain[5])) | (soc_ethmac_rx_cdc_graycounter0_q[4:0] != soc_ethmac_rx_cdc_consume_wdomain[4:0]));
assign soc_ethmac_rx_cdc_asyncfifo_readable = (soc_ethmac_rx_cdc_graycounter1_q != soc_ethmac_rx_cdc_produce_rdomain);
assign soc_ethmac_rx_cdc_wrport_adr = soc_ethmac_rx_cdc_graycounter0_q_binary[5:0];
assign soc_ethmac_rx_cdc_wrport_dat_w = soc_ethmac_rx_cdc_asyncfifo_din;
assign soc_ethmac_rx_cdc_wrport_we = soc_ethmac_rx_cdc_graycounter0_ce;
assign soc_ethmac_rx_cdc_rdport_adr = soc_ethmac_rx_cdc_graycounter1_q_next_binary[5:0];
assign soc_ethmac_rx_cdc_asyncfifo_dout = soc_ethmac_rx_cdc_rdport_dat_r;
always @(*) begin
	soc_ethmac_rx_cdc_graycounter0_q_next_binary <= 7'd0;
	if (soc_ethmac_rx_cdc_graycounter0_ce) begin
		soc_ethmac_rx_cdc_graycounter0_q_next_binary <= (soc_ethmac_rx_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		soc_ethmac_rx_cdc_graycounter0_q_next_binary <= soc_ethmac_rx_cdc_graycounter0_q_binary;
	end
end
assign soc_ethmac_rx_cdc_graycounter0_q_next = (soc_ethmac_rx_cdc_graycounter0_q_next_binary ^ soc_ethmac_rx_cdc_graycounter0_q_next_binary[6:1]);
always @(*) begin
	soc_ethmac_rx_cdc_graycounter1_q_next_binary <= 7'd0;
	if (soc_ethmac_rx_cdc_graycounter1_ce) begin
		soc_ethmac_rx_cdc_graycounter1_q_next_binary <= (soc_ethmac_rx_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		soc_ethmac_rx_cdc_graycounter1_q_next_binary <= soc_ethmac_rx_cdc_graycounter1_q_binary;
	end
end
assign soc_ethmac_rx_cdc_graycounter1_q_next = (soc_ethmac_rx_cdc_graycounter1_q_next_binary ^ soc_ethmac_rx_cdc_graycounter1_q_next_binary[6:1]);
assign soc_ethmac_tx_converter_sink_valid = soc_ethmac_tx_cdc_source_valid;
assign soc_ethmac_tx_cdc_source_ready = soc_ethmac_tx_converter_sink_ready;
assign soc_ethmac_tx_converter_sink_first = soc_ethmac_tx_cdc_source_first;
assign soc_ethmac_tx_converter_sink_last = soc_ethmac_tx_cdc_source_last;
assign soc_ethmac_tx_converter_sink_payload_data = soc_ethmac_tx_cdc_source_payload_data;
assign soc_ethmac_tx_converter_sink_payload_last_be = soc_ethmac_tx_cdc_source_payload_last_be;
assign soc_ethmac_tx_converter_sink_payload_error = soc_ethmac_tx_cdc_source_payload_error;
assign soc_ethmac_tx_last_be_sink_valid = soc_ethmac_tx_converter_source_valid;
assign soc_ethmac_tx_converter_source_ready = soc_ethmac_tx_last_be_sink_ready;
assign soc_ethmac_tx_last_be_sink_first = soc_ethmac_tx_converter_source_first;
assign soc_ethmac_tx_last_be_sink_last = soc_ethmac_tx_converter_source_last;
assign soc_ethmac_tx_last_be_sink_payload_data = soc_ethmac_tx_converter_source_payload_data;
assign soc_ethmac_tx_last_be_sink_payload_last_be = soc_ethmac_tx_converter_source_payload_last_be;
assign soc_ethmac_tx_last_be_sink_payload_error = soc_ethmac_tx_converter_source_payload_error;
assign soc_ethmac_padding_inserter_sink_valid = soc_ethmac_tx_last_be_source_valid;
assign soc_ethmac_tx_last_be_source_ready = soc_ethmac_padding_inserter_sink_ready;
assign soc_ethmac_padding_inserter_sink_first = soc_ethmac_tx_last_be_source_first;
assign soc_ethmac_padding_inserter_sink_last = soc_ethmac_tx_last_be_source_last;
assign soc_ethmac_padding_inserter_sink_payload_data = soc_ethmac_tx_last_be_source_payload_data;
assign soc_ethmac_padding_inserter_sink_payload_last_be = soc_ethmac_tx_last_be_source_payload_last_be;
assign soc_ethmac_padding_inserter_sink_payload_error = soc_ethmac_tx_last_be_source_payload_error;
assign soc_ethmac_crc32_inserter_sink_valid = soc_ethmac_padding_inserter_source_valid;
assign soc_ethmac_padding_inserter_source_ready = soc_ethmac_crc32_inserter_sink_ready;
assign soc_ethmac_crc32_inserter_sink_first = soc_ethmac_padding_inserter_source_first;
assign soc_ethmac_crc32_inserter_sink_last = soc_ethmac_padding_inserter_source_last;
assign soc_ethmac_crc32_inserter_sink_payload_data = soc_ethmac_padding_inserter_source_payload_data;
assign soc_ethmac_crc32_inserter_sink_payload_last_be = soc_ethmac_padding_inserter_source_payload_last_be;
assign soc_ethmac_crc32_inserter_sink_payload_error = soc_ethmac_padding_inserter_source_payload_error;
assign soc_ethmac_preamble_inserter_sink_valid = soc_ethmac_crc32_inserter_source_valid;
assign soc_ethmac_crc32_inserter_source_ready = soc_ethmac_preamble_inserter_sink_ready;
assign soc_ethmac_preamble_inserter_sink_first = soc_ethmac_crc32_inserter_source_first;
assign soc_ethmac_preamble_inserter_sink_last = soc_ethmac_crc32_inserter_source_last;
assign soc_ethmac_preamble_inserter_sink_payload_data = soc_ethmac_crc32_inserter_source_payload_data;
assign soc_ethmac_preamble_inserter_sink_payload_last_be = soc_ethmac_crc32_inserter_source_payload_last_be;
assign soc_ethmac_preamble_inserter_sink_payload_error = soc_ethmac_crc32_inserter_source_payload_error;
assign soc_ethmac_tx_gap_inserter_sink_valid = soc_ethmac_preamble_inserter_source_valid;
assign soc_ethmac_preamble_inserter_source_ready = soc_ethmac_tx_gap_inserter_sink_ready;
assign soc_ethmac_tx_gap_inserter_sink_first = soc_ethmac_preamble_inserter_source_first;
assign soc_ethmac_tx_gap_inserter_sink_last = soc_ethmac_preamble_inserter_source_last;
assign soc_ethmac_tx_gap_inserter_sink_payload_data = soc_ethmac_preamble_inserter_source_payload_data;
assign soc_ethmac_tx_gap_inserter_sink_payload_last_be = soc_ethmac_preamble_inserter_source_payload_last_be;
assign soc_ethmac_tx_gap_inserter_sink_payload_error = soc_ethmac_preamble_inserter_source_payload_error;
assign soc_ethphy_sink_valid = soc_ethmac_tx_gap_inserter_source_valid;
assign soc_ethmac_tx_gap_inserter_source_ready = soc_ethphy_sink_ready;
assign soc_ethphy_sink_first = soc_ethmac_tx_gap_inserter_source_first;
assign soc_ethphy_sink_last = soc_ethmac_tx_gap_inserter_source_last;
assign soc_ethphy_sink_payload_data = soc_ethmac_tx_gap_inserter_source_payload_data;
assign soc_ethphy_sink_payload_last_be = soc_ethmac_tx_gap_inserter_source_payload_last_be;
assign soc_ethphy_sink_payload_error = soc_ethmac_tx_gap_inserter_source_payload_error;
assign soc_ethmac_rx_gap_checker_sink_valid = soc_ethphy_source_valid;
assign soc_ethphy_source_ready = soc_ethmac_rx_gap_checker_sink_ready;
assign soc_ethmac_rx_gap_checker_sink_first = soc_ethphy_source_first;
assign soc_ethmac_rx_gap_checker_sink_last = soc_ethphy_source_last;
assign soc_ethmac_rx_gap_checker_sink_payload_data = soc_ethphy_source_payload_data;
assign soc_ethmac_rx_gap_checker_sink_payload_last_be = soc_ethphy_source_payload_last_be;
assign soc_ethmac_rx_gap_checker_sink_payload_error = soc_ethphy_source_payload_error;
assign soc_ethmac_preamble_checker_sink_valid = soc_ethmac_rx_gap_checker_source_valid;
assign soc_ethmac_rx_gap_checker_source_ready = soc_ethmac_preamble_checker_sink_ready;
assign soc_ethmac_preamble_checker_sink_first = soc_ethmac_rx_gap_checker_source_first;
assign soc_ethmac_preamble_checker_sink_last = soc_ethmac_rx_gap_checker_source_last;
assign soc_ethmac_preamble_checker_sink_payload_data = soc_ethmac_rx_gap_checker_source_payload_data;
assign soc_ethmac_preamble_checker_sink_payload_last_be = soc_ethmac_rx_gap_checker_source_payload_last_be;
assign soc_ethmac_preamble_checker_sink_payload_error = soc_ethmac_rx_gap_checker_source_payload_error;
assign soc_ethmac_crc32_checker_sink_sink_valid = soc_ethmac_preamble_checker_source_valid;
assign soc_ethmac_preamble_checker_source_ready = soc_ethmac_crc32_checker_sink_sink_ready;
assign soc_ethmac_crc32_checker_sink_sink_first = soc_ethmac_preamble_checker_source_first;
assign soc_ethmac_crc32_checker_sink_sink_last = soc_ethmac_preamble_checker_source_last;
assign soc_ethmac_crc32_checker_sink_sink_payload_data = soc_ethmac_preamble_checker_source_payload_data;
assign soc_ethmac_crc32_checker_sink_sink_payload_last_be = soc_ethmac_preamble_checker_source_payload_last_be;
assign soc_ethmac_crc32_checker_sink_sink_payload_error = soc_ethmac_preamble_checker_source_payload_error;
assign soc_ethmac_padding_checker_sink_valid = soc_ethmac_crc32_checker_source_source_valid;
assign soc_ethmac_crc32_checker_source_source_ready = soc_ethmac_padding_checker_sink_ready;
assign soc_ethmac_padding_checker_sink_first = soc_ethmac_crc32_checker_source_source_first;
assign soc_ethmac_padding_checker_sink_last = soc_ethmac_crc32_checker_source_source_last;
assign soc_ethmac_padding_checker_sink_payload_data = soc_ethmac_crc32_checker_source_source_payload_data;
assign soc_ethmac_padding_checker_sink_payload_last_be = soc_ethmac_crc32_checker_source_source_payload_last_be;
assign soc_ethmac_padding_checker_sink_payload_error = soc_ethmac_crc32_checker_source_source_payload_error;
assign soc_ethmac_rx_last_be_sink_valid = soc_ethmac_padding_checker_source_valid;
assign soc_ethmac_padding_checker_source_ready = soc_ethmac_rx_last_be_sink_ready;
assign soc_ethmac_rx_last_be_sink_first = soc_ethmac_padding_checker_source_first;
assign soc_ethmac_rx_last_be_sink_last = soc_ethmac_padding_checker_source_last;
assign soc_ethmac_rx_last_be_sink_payload_data = soc_ethmac_padding_checker_source_payload_data;
assign soc_ethmac_rx_last_be_sink_payload_last_be = soc_ethmac_padding_checker_source_payload_last_be;
assign soc_ethmac_rx_last_be_sink_payload_error = soc_ethmac_padding_checker_source_payload_error;
assign soc_ethmac_rx_converter_sink_valid = soc_ethmac_rx_last_be_source_valid;
assign soc_ethmac_rx_last_be_source_ready = soc_ethmac_rx_converter_sink_ready;
assign soc_ethmac_rx_converter_sink_first = soc_ethmac_rx_last_be_source_first;
assign soc_ethmac_rx_converter_sink_last = soc_ethmac_rx_last_be_source_last;
assign soc_ethmac_rx_converter_sink_payload_data = soc_ethmac_rx_last_be_source_payload_data;
assign soc_ethmac_rx_converter_sink_payload_last_be = soc_ethmac_rx_last_be_source_payload_last_be;
assign soc_ethmac_rx_converter_sink_payload_error = soc_ethmac_rx_last_be_source_payload_error;
assign soc_ethmac_rx_cdc_sink_valid = soc_ethmac_rx_converter_source_valid;
assign soc_ethmac_rx_converter_source_ready = soc_ethmac_rx_cdc_sink_ready;
assign soc_ethmac_rx_cdc_sink_first = soc_ethmac_rx_converter_source_first;
assign soc_ethmac_rx_cdc_sink_last = soc_ethmac_rx_converter_source_last;
assign soc_ethmac_rx_cdc_sink_payload_data = soc_ethmac_rx_converter_source_payload_data;
assign soc_ethmac_rx_cdc_sink_payload_last_be = soc_ethmac_rx_converter_source_payload_last_be;
assign soc_ethmac_rx_cdc_sink_payload_error = soc_ethmac_rx_converter_source_payload_error;
assign soc_ethmac_writer_sink_sink_valid = soc_ethmac_sink_valid;
assign soc_ethmac_sink_ready = soc_ethmac_writer_sink_sink_ready;
assign soc_ethmac_writer_sink_sink_first = soc_ethmac_sink_first;
assign soc_ethmac_writer_sink_sink_last = soc_ethmac_sink_last;
assign soc_ethmac_writer_sink_sink_payload_data = soc_ethmac_sink_payload_data;
assign soc_ethmac_writer_sink_sink_payload_last_be = soc_ethmac_sink_payload_last_be;
assign soc_ethmac_writer_sink_sink_payload_error = soc_ethmac_sink_payload_error;
assign soc_ethmac_source_valid = soc_ethmac_reader_source_source_valid;
assign soc_ethmac_reader_source_source_ready = soc_ethmac_source_ready;
assign soc_ethmac_source_first = soc_ethmac_reader_source_source_first;
assign soc_ethmac_source_last = soc_ethmac_reader_source_source_last;
assign soc_ethmac_source_payload_data = soc_ethmac_reader_source_source_payload_data;
assign soc_ethmac_source_payload_last_be = soc_ethmac_reader_source_source_payload_last_be;
assign soc_ethmac_source_payload_error = soc_ethmac_reader_source_source_payload_error;
always @(*) begin
	soc_ethmac_writer_increment <= 3'd0;
	if (soc_ethmac_writer_sink_sink_payload_last_be[3]) begin
		soc_ethmac_writer_increment <= 1'd1;
	end else begin
		if (soc_ethmac_writer_sink_sink_payload_last_be[2]) begin
			soc_ethmac_writer_increment <= 2'd2;
		end else begin
			if (soc_ethmac_writer_sink_sink_payload_last_be[1]) begin
				soc_ethmac_writer_increment <= 2'd3;
			end else begin
				soc_ethmac_writer_increment <= 3'd4;
			end
		end
	end
end
assign soc_ethmac_writer_fifo_sink_payload_slot = soc_ethmac_writer_slot;
assign soc_ethmac_writer_fifo_sink_payload_length = soc_ethmac_writer_counter;
assign soc_ethmac_writer_fifo_source_ready = soc_ethmac_writer_available_clear;
assign soc_ethmac_writer_available_trigger = soc_ethmac_writer_fifo_source_valid;
assign soc_ethmac_writer_slot_status = soc_ethmac_writer_fifo_source_payload_slot;
assign soc_ethmac_writer_length_status = soc_ethmac_writer_fifo_source_payload_length;
always @(*) begin
	soc_ethmac_writer_memory0_we <= 1'd0;
	soc_ethmac_writer_memory0_dat_w <= 32'd0;
	soc_ethmac_writer_memory1_adr <= 9'd0;
	soc_ethmac_writer_memory1_we <= 1'd0;
	soc_ethmac_writer_memory0_adr <= 9'd0;
	soc_ethmac_writer_memory1_dat_w <= 32'd0;
	case (soc_ethmac_writer_slot)
		1'd0: begin
			soc_ethmac_writer_memory0_adr <= soc_ethmac_writer_counter[31:2];
			soc_ethmac_writer_memory0_dat_w <= soc_ethmac_writer_sink_sink_payload_data;
			if ((soc_ethmac_writer_sink_sink_valid & soc_ethmac_writer_ongoing)) begin
				soc_ethmac_writer_memory0_we <= 4'd15;
			end
		end
		1'd1: begin
			soc_ethmac_writer_memory1_adr <= soc_ethmac_writer_counter[31:2];
			soc_ethmac_writer_memory1_dat_w <= soc_ethmac_writer_sink_sink_payload_data;
			if ((soc_ethmac_writer_sink_sink_valid & soc_ethmac_writer_ongoing)) begin
				soc_ethmac_writer_memory1_we <= 4'd15;
			end
		end
	endcase
end
assign soc_ethmac_writer_status_w = soc_ethmac_writer_available_status;
always @(*) begin
	soc_ethmac_writer_available_clear <= 1'd0;
	if ((soc_ethmac_writer_pending_re & soc_ethmac_writer_pending_r)) begin
		soc_ethmac_writer_available_clear <= 1'd1;
	end
end
assign soc_ethmac_writer_pending_w = soc_ethmac_writer_available_pending;
assign soc_ethmac_writer_irq = (soc_ethmac_writer_pending_w & soc_ethmac_writer_storage);
assign soc_ethmac_writer_available_status = soc_ethmac_writer_available_trigger;
assign soc_ethmac_writer_available_pending = soc_ethmac_writer_available_trigger;
assign soc_ethmac_writer_fifo_syncfifo_din = {soc_ethmac_writer_fifo_fifo_in_last, soc_ethmac_writer_fifo_fifo_in_first, soc_ethmac_writer_fifo_fifo_in_payload_length, soc_ethmac_writer_fifo_fifo_in_payload_slot};
assign {soc_ethmac_writer_fifo_fifo_out_last, soc_ethmac_writer_fifo_fifo_out_first, soc_ethmac_writer_fifo_fifo_out_payload_length, soc_ethmac_writer_fifo_fifo_out_payload_slot} = soc_ethmac_writer_fifo_syncfifo_dout;
assign soc_ethmac_writer_fifo_sink_ready = soc_ethmac_writer_fifo_syncfifo_writable;
assign soc_ethmac_writer_fifo_syncfifo_we = soc_ethmac_writer_fifo_sink_valid;
assign soc_ethmac_writer_fifo_fifo_in_first = soc_ethmac_writer_fifo_sink_first;
assign soc_ethmac_writer_fifo_fifo_in_last = soc_ethmac_writer_fifo_sink_last;
assign soc_ethmac_writer_fifo_fifo_in_payload_slot = soc_ethmac_writer_fifo_sink_payload_slot;
assign soc_ethmac_writer_fifo_fifo_in_payload_length = soc_ethmac_writer_fifo_sink_payload_length;
assign soc_ethmac_writer_fifo_source_valid = soc_ethmac_writer_fifo_syncfifo_readable;
assign soc_ethmac_writer_fifo_source_first = soc_ethmac_writer_fifo_fifo_out_first;
assign soc_ethmac_writer_fifo_source_last = soc_ethmac_writer_fifo_fifo_out_last;
assign soc_ethmac_writer_fifo_source_payload_slot = soc_ethmac_writer_fifo_fifo_out_payload_slot;
assign soc_ethmac_writer_fifo_source_payload_length = soc_ethmac_writer_fifo_fifo_out_payload_length;
assign soc_ethmac_writer_fifo_syncfifo_re = soc_ethmac_writer_fifo_source_ready;
always @(*) begin
	soc_ethmac_writer_fifo_wrport_adr <= 1'd0;
	if (soc_ethmac_writer_fifo_replace) begin
		soc_ethmac_writer_fifo_wrport_adr <= (soc_ethmac_writer_fifo_produce - 1'd1);
	end else begin
		soc_ethmac_writer_fifo_wrport_adr <= soc_ethmac_writer_fifo_produce;
	end
end
assign soc_ethmac_writer_fifo_wrport_dat_w = soc_ethmac_writer_fifo_syncfifo_din;
assign soc_ethmac_writer_fifo_wrport_we = (soc_ethmac_writer_fifo_syncfifo_we & (soc_ethmac_writer_fifo_syncfifo_writable | soc_ethmac_writer_fifo_replace));
assign soc_ethmac_writer_fifo_do_read = (soc_ethmac_writer_fifo_syncfifo_readable & soc_ethmac_writer_fifo_syncfifo_re);
assign soc_ethmac_writer_fifo_rdport_adr = soc_ethmac_writer_fifo_consume;
assign soc_ethmac_writer_fifo_syncfifo_dout = soc_ethmac_writer_fifo_rdport_dat_r;
assign soc_ethmac_writer_fifo_syncfifo_writable = (soc_ethmac_writer_fifo_level != 2'd2);
assign soc_ethmac_writer_fifo_syncfifo_readable = (soc_ethmac_writer_fifo_level != 1'd0);
always @(*) begin
	soc_ethmac_writer_slot_ce <= 1'd0;
	vns_liteethmacsramwriter_next_state <= 2'd0;
	soc_ethmac_writer_ongoing <= 1'd0;
	soc_ethmac_writer_fifo_sink_valid <= 1'd0;
	soc_ethmac_writer_counter_reset <= 1'd0;
	soc_ethmac_writer_counter_ce <= 1'd0;
	vns_liteethmacsramwriter_next_state <= vns_liteethmacsramwriter_state;
	case (vns_liteethmacsramwriter_state)
		1'd1: begin
			soc_ethmac_writer_counter_ce <= soc_ethmac_writer_sink_sink_valid;
			soc_ethmac_writer_ongoing <= (soc_ethmac_writer_counter < 11'd1530);
			if ((soc_ethmac_writer_sink_sink_valid & soc_ethmac_writer_sink_sink_last)) begin
				if (((soc_ethmac_writer_sink_sink_payload_error & soc_ethmac_writer_sink_sink_payload_last_be) != 1'd0)) begin
					vns_liteethmacsramwriter_next_state <= 2'd2;
				end else begin
					vns_liteethmacsramwriter_next_state <= 2'd3;
				end
			end
		end
		2'd2: begin
			soc_ethmac_writer_counter_reset <= 1'd1;
			vns_liteethmacsramwriter_next_state <= 1'd0;
		end
		2'd3: begin
			soc_ethmac_writer_counter_reset <= 1'd1;
			soc_ethmac_writer_slot_ce <= 1'd1;
			soc_ethmac_writer_fifo_sink_valid <= 1'd1;
			vns_liteethmacsramwriter_next_state <= 1'd0;
		end
		default: begin
			if (soc_ethmac_writer_sink_sink_valid) begin
				if (soc_ethmac_writer_fifo_sink_ready) begin
					soc_ethmac_writer_ongoing <= 1'd1;
					soc_ethmac_writer_counter_ce <= 1'd1;
					vns_liteethmacsramwriter_next_state <= 1'd1;
				end
			end
		end
	endcase
end
assign soc_ethmac_reader_fifo_sink_valid = soc_ethmac_reader_start_re;
assign soc_ethmac_reader_fifo_sink_payload_slot = soc_ethmac_reader_slot_storage;
assign soc_ethmac_reader_fifo_sink_payload_length = soc_ethmac_reader_length_storage;
assign soc_ethmac_reader_ready_status = soc_ethmac_reader_fifo_sink_ready;
always @(*) begin
	soc_ethmac_reader_source_source_payload_last_be <= 4'd0;
	if (soc_ethmac_reader_last) begin
		if ((soc_ethmac_reader_fifo_source_payload_length[1:0] == 2'd3)) begin
			soc_ethmac_reader_source_source_payload_last_be <= 2'd2;
		end else begin
			if ((soc_ethmac_reader_fifo_source_payload_length[1:0] == 2'd2)) begin
				soc_ethmac_reader_source_source_payload_last_be <= 3'd4;
			end else begin
				if ((soc_ethmac_reader_fifo_source_payload_length[1:0] == 1'd1)) begin
					soc_ethmac_reader_source_source_payload_last_be <= 4'd8;
				end else begin
					soc_ethmac_reader_source_source_payload_last_be <= 1'd1;
				end
			end
		end
	end
end
assign soc_ethmac_reader_last = (soc_ethmac_reader_counter >= soc_ethmac_reader_fifo_source_payload_length);
assign soc_ethmac_reader_memory0_adr = soc_ethmac_reader_counter[10:2];
assign soc_ethmac_reader_memory1_adr = soc_ethmac_reader_counter[10:2];
always @(*) begin
	soc_ethmac_reader_source_source_payload_data <= 32'd0;
	case (soc_ethmac_reader_fifo_source_payload_slot)
		1'd0: begin
			soc_ethmac_reader_source_source_payload_data <= soc_ethmac_reader_memory0_dat_r;
		end
		1'd1: begin
			soc_ethmac_reader_source_source_payload_data <= soc_ethmac_reader_memory1_dat_r;
		end
	endcase
end
assign soc_ethmac_reader_eventmanager_status_w = soc_ethmac_reader_done_status;
always @(*) begin
	soc_ethmac_reader_done_clear <= 1'd0;
	if ((soc_ethmac_reader_eventmanager_pending_re & soc_ethmac_reader_eventmanager_pending_r)) begin
		soc_ethmac_reader_done_clear <= 1'd1;
	end
end
assign soc_ethmac_reader_eventmanager_pending_w = soc_ethmac_reader_done_pending;
assign soc_ethmac_reader_irq = (soc_ethmac_reader_eventmanager_pending_w & soc_ethmac_reader_eventmanager_storage);
assign soc_ethmac_reader_done_status = 1'd0;
assign soc_ethmac_reader_fifo_syncfifo_din = {soc_ethmac_reader_fifo_fifo_in_last, soc_ethmac_reader_fifo_fifo_in_first, soc_ethmac_reader_fifo_fifo_in_payload_length, soc_ethmac_reader_fifo_fifo_in_payload_slot};
assign {soc_ethmac_reader_fifo_fifo_out_last, soc_ethmac_reader_fifo_fifo_out_first, soc_ethmac_reader_fifo_fifo_out_payload_length, soc_ethmac_reader_fifo_fifo_out_payload_slot} = soc_ethmac_reader_fifo_syncfifo_dout;
assign soc_ethmac_reader_fifo_sink_ready = soc_ethmac_reader_fifo_syncfifo_writable;
assign soc_ethmac_reader_fifo_syncfifo_we = soc_ethmac_reader_fifo_sink_valid;
assign soc_ethmac_reader_fifo_fifo_in_first = soc_ethmac_reader_fifo_sink_first;
assign soc_ethmac_reader_fifo_fifo_in_last = soc_ethmac_reader_fifo_sink_last;
assign soc_ethmac_reader_fifo_fifo_in_payload_slot = soc_ethmac_reader_fifo_sink_payload_slot;
assign soc_ethmac_reader_fifo_fifo_in_payload_length = soc_ethmac_reader_fifo_sink_payload_length;
assign soc_ethmac_reader_fifo_source_valid = soc_ethmac_reader_fifo_syncfifo_readable;
assign soc_ethmac_reader_fifo_source_first = soc_ethmac_reader_fifo_fifo_out_first;
assign soc_ethmac_reader_fifo_source_last = soc_ethmac_reader_fifo_fifo_out_last;
assign soc_ethmac_reader_fifo_source_payload_slot = soc_ethmac_reader_fifo_fifo_out_payload_slot;
assign soc_ethmac_reader_fifo_source_payload_length = soc_ethmac_reader_fifo_fifo_out_payload_length;
assign soc_ethmac_reader_fifo_syncfifo_re = soc_ethmac_reader_fifo_source_ready;
always @(*) begin
	soc_ethmac_reader_fifo_wrport_adr <= 1'd0;
	if (soc_ethmac_reader_fifo_replace) begin
		soc_ethmac_reader_fifo_wrport_adr <= (soc_ethmac_reader_fifo_produce - 1'd1);
	end else begin
		soc_ethmac_reader_fifo_wrport_adr <= soc_ethmac_reader_fifo_produce;
	end
end
assign soc_ethmac_reader_fifo_wrport_dat_w = soc_ethmac_reader_fifo_syncfifo_din;
assign soc_ethmac_reader_fifo_wrport_we = (soc_ethmac_reader_fifo_syncfifo_we & (soc_ethmac_reader_fifo_syncfifo_writable | soc_ethmac_reader_fifo_replace));
assign soc_ethmac_reader_fifo_do_read = (soc_ethmac_reader_fifo_syncfifo_readable & soc_ethmac_reader_fifo_syncfifo_re);
assign soc_ethmac_reader_fifo_rdport_adr = soc_ethmac_reader_fifo_consume;
assign soc_ethmac_reader_fifo_syncfifo_dout = soc_ethmac_reader_fifo_rdport_dat_r;
assign soc_ethmac_reader_fifo_syncfifo_writable = (soc_ethmac_reader_fifo_level != 2'd2);
assign soc_ethmac_reader_fifo_syncfifo_readable = (soc_ethmac_reader_fifo_level != 1'd0);
always @(*) begin
	soc_ethmac_reader_source_source_last <= 1'd0;
	soc_ethmac_reader_done_trigger <= 1'd0;
	vns_liteethmacsramreader_next_state <= 2'd0;
	soc_ethmac_reader_counter_reset <= 1'd0;
	soc_ethmac_reader_source_source_valid <= 1'd0;
	soc_ethmac_reader_counter_ce <= 1'd0;
	soc_ethmac_reader_fifo_source_ready <= 1'd0;
	vns_liteethmacsramreader_next_state <= vns_liteethmacsramreader_state;
	case (vns_liteethmacsramreader_state)
		1'd1: begin
			soc_ethmac_reader_source_source_valid <= 1'd1;
			soc_ethmac_reader_source_source_last <= soc_ethmac_reader_last;
			if (soc_ethmac_reader_source_source_ready) begin
				soc_ethmac_reader_counter_ce <= 1'd1;
				if (soc_ethmac_reader_last) begin
					vns_liteethmacsramreader_next_state <= 2'd2;
				end
			end
		end
		2'd2: begin
			soc_ethmac_reader_fifo_source_ready <= 1'd1;
			soc_ethmac_reader_done_trigger <= 1'd1;
			soc_ethmac_reader_counter_reset <= 1'd1;
			vns_liteethmacsramreader_next_state <= 1'd0;
		end
		default: begin
			if (soc_ethmac_reader_fifo_source_valid) begin
				soc_ethmac_reader_counter_ce <= 1'd1;
				vns_liteethmacsramreader_next_state <= 1'd1;
			end
		end
	endcase
end
assign soc_ethmac_ev_irq = (soc_ethmac_writer_irq | soc_ethmac_reader_irq);
assign soc_ethmac_sram0_adr0 = soc_ethmac_sram0_bus_adr0[8:0];
assign soc_ethmac_sram0_bus_dat_r0 = soc_ethmac_sram0_dat_r0;
assign soc_ethmac_sram1_adr0 = soc_ethmac_sram1_bus_adr0[8:0];
assign soc_ethmac_sram1_bus_dat_r0 = soc_ethmac_sram1_dat_r0;
always @(*) begin
	soc_ethmac_sram0_we <= 4'd0;
	soc_ethmac_sram0_we[0] <= (((soc_ethmac_sram0_bus_cyc1 & soc_ethmac_sram0_bus_stb1) & soc_ethmac_sram0_bus_we1) & soc_ethmac_sram0_bus_sel1[0]);
	soc_ethmac_sram0_we[1] <= (((soc_ethmac_sram0_bus_cyc1 & soc_ethmac_sram0_bus_stb1) & soc_ethmac_sram0_bus_we1) & soc_ethmac_sram0_bus_sel1[1]);
	soc_ethmac_sram0_we[2] <= (((soc_ethmac_sram0_bus_cyc1 & soc_ethmac_sram0_bus_stb1) & soc_ethmac_sram0_bus_we1) & soc_ethmac_sram0_bus_sel1[2]);
	soc_ethmac_sram0_we[3] <= (((soc_ethmac_sram0_bus_cyc1 & soc_ethmac_sram0_bus_stb1) & soc_ethmac_sram0_bus_we1) & soc_ethmac_sram0_bus_sel1[3]);
end
assign soc_ethmac_sram0_adr1 = soc_ethmac_sram0_bus_adr1[8:0];
assign soc_ethmac_sram0_bus_dat_r1 = soc_ethmac_sram0_dat_r1;
assign soc_ethmac_sram0_dat_w = soc_ethmac_sram0_bus_dat_w1;
always @(*) begin
	soc_ethmac_sram1_we <= 4'd0;
	soc_ethmac_sram1_we[0] <= (((soc_ethmac_sram1_bus_cyc1 & soc_ethmac_sram1_bus_stb1) & soc_ethmac_sram1_bus_we1) & soc_ethmac_sram1_bus_sel1[0]);
	soc_ethmac_sram1_we[1] <= (((soc_ethmac_sram1_bus_cyc1 & soc_ethmac_sram1_bus_stb1) & soc_ethmac_sram1_bus_we1) & soc_ethmac_sram1_bus_sel1[1]);
	soc_ethmac_sram1_we[2] <= (((soc_ethmac_sram1_bus_cyc1 & soc_ethmac_sram1_bus_stb1) & soc_ethmac_sram1_bus_we1) & soc_ethmac_sram1_bus_sel1[2]);
	soc_ethmac_sram1_we[3] <= (((soc_ethmac_sram1_bus_cyc1 & soc_ethmac_sram1_bus_stb1) & soc_ethmac_sram1_bus_we1) & soc_ethmac_sram1_bus_sel1[3]);
end
assign soc_ethmac_sram1_adr1 = soc_ethmac_sram1_bus_adr1[8:0];
assign soc_ethmac_sram1_bus_dat_r1 = soc_ethmac_sram1_dat_r1;
assign soc_ethmac_sram1_dat_w = soc_ethmac_sram1_bus_dat_w1;
always @(*) begin
	soc_ethmac_slave_sel <= 4'd0;
	soc_ethmac_slave_sel[0] <= (soc_ethmac_bus_adr[10:9] == 1'd0);
	soc_ethmac_slave_sel[1] <= (soc_ethmac_bus_adr[10:9] == 1'd1);
	soc_ethmac_slave_sel[2] <= (soc_ethmac_bus_adr[10:9] == 2'd2);
	soc_ethmac_slave_sel[3] <= (soc_ethmac_bus_adr[10:9] == 2'd3);
end
assign soc_ethmac_sram0_bus_adr0 = soc_ethmac_bus_adr;
assign soc_ethmac_sram0_bus_dat_w0 = soc_ethmac_bus_dat_w;
assign soc_ethmac_sram0_bus_sel0 = soc_ethmac_bus_sel;
assign soc_ethmac_sram0_bus_stb0 = soc_ethmac_bus_stb;
assign soc_ethmac_sram0_bus_we0 = soc_ethmac_bus_we;
assign soc_ethmac_sram0_bus_cti0 = soc_ethmac_bus_cti;
assign soc_ethmac_sram0_bus_bte0 = soc_ethmac_bus_bte;
assign soc_ethmac_sram1_bus_adr0 = soc_ethmac_bus_adr;
assign soc_ethmac_sram1_bus_dat_w0 = soc_ethmac_bus_dat_w;
assign soc_ethmac_sram1_bus_sel0 = soc_ethmac_bus_sel;
assign soc_ethmac_sram1_bus_stb0 = soc_ethmac_bus_stb;
assign soc_ethmac_sram1_bus_we0 = soc_ethmac_bus_we;
assign soc_ethmac_sram1_bus_cti0 = soc_ethmac_bus_cti;
assign soc_ethmac_sram1_bus_bte0 = soc_ethmac_bus_bte;
assign soc_ethmac_sram0_bus_adr1 = soc_ethmac_bus_adr;
assign soc_ethmac_sram0_bus_dat_w1 = soc_ethmac_bus_dat_w;
assign soc_ethmac_sram0_bus_sel1 = soc_ethmac_bus_sel;
assign soc_ethmac_sram0_bus_stb1 = soc_ethmac_bus_stb;
assign soc_ethmac_sram0_bus_we1 = soc_ethmac_bus_we;
assign soc_ethmac_sram0_bus_cti1 = soc_ethmac_bus_cti;
assign soc_ethmac_sram0_bus_bte1 = soc_ethmac_bus_bte;
assign soc_ethmac_sram1_bus_adr1 = soc_ethmac_bus_adr;
assign soc_ethmac_sram1_bus_dat_w1 = soc_ethmac_bus_dat_w;
assign soc_ethmac_sram1_bus_sel1 = soc_ethmac_bus_sel;
assign soc_ethmac_sram1_bus_stb1 = soc_ethmac_bus_stb;
assign soc_ethmac_sram1_bus_we1 = soc_ethmac_bus_we;
assign soc_ethmac_sram1_bus_cti1 = soc_ethmac_bus_cti;
assign soc_ethmac_sram1_bus_bte1 = soc_ethmac_bus_bte;
assign soc_ethmac_sram0_bus_cyc0 = (soc_ethmac_bus_cyc & soc_ethmac_slave_sel[0]);
assign soc_ethmac_sram1_bus_cyc0 = (soc_ethmac_bus_cyc & soc_ethmac_slave_sel[1]);
assign soc_ethmac_sram0_bus_cyc1 = (soc_ethmac_bus_cyc & soc_ethmac_slave_sel[2]);
assign soc_ethmac_sram1_bus_cyc1 = (soc_ethmac_bus_cyc & soc_ethmac_slave_sel[3]);
assign soc_ethmac_bus_ack = (((soc_ethmac_sram0_bus_ack0 | soc_ethmac_sram1_bus_ack0) | soc_ethmac_sram0_bus_ack1) | soc_ethmac_sram1_bus_ack1);
assign soc_ethmac_bus_err = (((soc_ethmac_sram0_bus_err0 | soc_ethmac_sram1_bus_err0) | soc_ethmac_sram0_bus_err1) | soc_ethmac_sram1_bus_err1);
assign soc_ethmac_bus_dat_r = (((({32{soc_ethmac_slave_sel_r[0]}} & soc_ethmac_sram0_bus_dat_r0) | ({32{soc_ethmac_slave_sel_r[1]}} & soc_ethmac_sram1_bus_dat_r0)) | ({32{soc_ethmac_slave_sel_r[2]}} & soc_ethmac_sram0_bus_dat_r1)) | ({32{soc_ethmac_slave_sel_r[3]}} & soc_ethmac_sram1_bus_dat_r1));
assign soc_charsync0_raw_data = soc_s7datacapture0_d;
assign soc_wer0_data = soc_charsync0_data;
assign soc_decoding0_valid_i = soc_charsync0_synced;
assign soc_decoding0_input = soc_charsync0_data;
assign soc_charsync1_raw_data = soc_s7datacapture1_d;
assign soc_wer1_data = soc_charsync1_data;
assign soc_decoding1_valid_i = soc_charsync1_synced;
assign soc_decoding1_input = soc_charsync1_data;
assign soc_charsync2_raw_data = soc_s7datacapture2_d;
assign soc_wer2_data = soc_charsync2_data;
assign soc_decoding2_valid_i = soc_charsync2_synced;
assign soc_decoding2_input = soc_charsync2_data;
assign soc_chansync_valid_i = ((soc_decoding0_valid_o & soc_decoding1_valid_o) & soc_decoding2_valid_o);
assign soc_chansync_data_in0_d = soc_decoding0_output_d;
assign soc_chansync_data_in0_c = soc_decoding0_output_c;
assign soc_chansync_data_in0_de = soc_decoding0_output_de;
assign soc_chansync_data_in1_d = soc_decoding1_output_d;
assign soc_chansync_data_in1_c = soc_decoding1_output_c;
assign soc_chansync_data_in1_de = soc_decoding1_output_de;
assign soc_chansync_data_in2_d = soc_decoding2_output_d;
assign soc_chansync_data_in2_c = soc_decoding2_output_c;
assign soc_chansync_data_in2_de = soc_decoding2_output_de;
assign soc_syncpol_valid_i = soc_chansync_chan_synced;
assign soc_syncpol_data_in0_d = soc_chansync_data_out0_d;
assign soc_syncpol_data_in0_c = soc_chansync_data_out0_c;
assign soc_syncpol_data_in0_de = soc_chansync_data_out0_de;
assign soc_syncpol_data_in1_d = soc_chansync_data_out1_d;
assign soc_syncpol_data_in1_c = soc_chansync_data_out1_c;
assign soc_syncpol_data_in1_de = soc_chansync_data_out1_de;
assign soc_syncpol_data_in2_d = soc_chansync_data_out2_d;
assign soc_syncpol_data_in2_c = soc_chansync_data_out2_c;
assign soc_syncpol_data_in2_de = soc_chansync_data_out2_de;
assign soc_resdetection_valid_i = soc_syncpol_valid_o;
assign soc_resdetection_de = soc_syncpol_de;
assign soc_resdetection_vsync = soc_syncpol_vsync;
assign soc_frame_valid_i = soc_syncpol_valid_o;
assign soc_frame_de = soc_syncpol_de;
assign soc_frame_vsync = soc_syncpol_vsync;
assign soc_frame_r = soc_syncpol_r;
assign soc_frame_g = soc_syncpol_g;
assign soc_frame_b = soc_syncpol_b;
assign soc_dma_frame_valid = soc_frame_frame_valid;
assign soc_frame_frame_ready = soc_dma_frame_ready;
assign soc_dma_frame_first = soc_frame_frame_first;
assign soc_dma_frame_last = soc_frame_frame_last;
assign soc_dma_frame_payload_sof = soc_frame_frame_payload_sof;
assign soc_dma_frame_payload_pixels = soc_frame_frame_payload_pixels;
assign soc_edid_status = 1'd1;
assign hdmi_in_hpd_en = soc_edid_storage;
assign soc_edid_sda_o = (~soc_edid_sda_drv_reg);
assign soc_edid_scl_rising = (soc_edid_scl_i & (~soc_edid_scl_r));
assign soc_edid_sda_rising = (soc_edid_sda_i & (~soc_edid_sda_r));
assign soc_edid_sda_falling = ((~soc_edid_sda_i) & soc_edid_sda_r);
assign soc_edid_start = (soc_edid_scl_i & soc_edid_sda_falling);
assign soc_edid_adr = soc_edid_offset_counter;
always @(*) begin
	soc_edid_sda_drv <= 1'd0;
	if (soc_edid_zero_drv) begin
		soc_edid_sda_drv <= 1'd1;
	end else begin
		if (soc_edid_data_drv) begin
			soc_edid_sda_drv <= (~soc_edid_data_bit);
		end
	end
end
always @(*) begin
	soc_edid_zero_drv <= 1'd0;
	soc_edid_oc_load <= 1'd0;
	soc_edid_oc_inc <= 1'd0;
	soc_edid_data_drv_en <= 1'd0;
	soc_edid_data_drv_stop <= 1'd0;
	vns_edid_next_state <= 4'd0;
	soc_edid_update_is_read <= 1'd0;
	vns_edid_next_state <= vns_edid_state;
	case (vns_edid_state)
		1'd1: begin
			if ((soc_edid_counter == 4'd8)) begin
				if ((soc_edid_din[7:1] == 7'd80)) begin
					soc_edid_update_is_read <= 1'd1;
					vns_edid_next_state <= 2'd2;
				end else begin
					vns_edid_next_state <= 1'd0;
				end
			end
			if (soc_edid_start) begin
				vns_edid_next_state <= 1'd1;
			end
			if ((~soc_edid_storage)) begin
				vns_edid_next_state <= 1'd0;
			end
		end
		2'd2: begin
			if ((~soc_edid_scl_i)) begin
				vns_edid_next_state <= 2'd3;
			end
			if (soc_edid_start) begin
				vns_edid_next_state <= 1'd1;
			end
			if ((~soc_edid_storage)) begin
				vns_edid_next_state <= 1'd0;
			end
		end
		2'd3: begin
			soc_edid_zero_drv <= 1'd1;
			if (soc_edid_scl_i) begin
				vns_edid_next_state <= 3'd4;
			end
			if (soc_edid_start) begin
				vns_edid_next_state <= 1'd1;
			end
			if ((~soc_edid_storage)) begin
				vns_edid_next_state <= 1'd0;
			end
		end
		3'd4: begin
			soc_edid_zero_drv <= 1'd1;
			if ((~soc_edid_scl_i)) begin
				if (soc_edid_is_read) begin
					vns_edid_next_state <= 4'd9;
				end else begin
					vns_edid_next_state <= 3'd5;
				end
			end
			if (soc_edid_start) begin
				vns_edid_next_state <= 1'd1;
			end
			if ((~soc_edid_storage)) begin
				vns_edid_next_state <= 1'd0;
			end
		end
		3'd5: begin
			if ((soc_edid_counter == 4'd8)) begin
				soc_edid_oc_load <= 1'd1;
				vns_edid_next_state <= 3'd6;
			end
			if (soc_edid_start) begin
				vns_edid_next_state <= 1'd1;
			end
			if ((~soc_edid_storage)) begin
				vns_edid_next_state <= 1'd0;
			end
		end
		3'd6: begin
			if ((~soc_edid_scl_i)) begin
				vns_edid_next_state <= 3'd7;
			end
			if (soc_edid_start) begin
				vns_edid_next_state <= 1'd1;
			end
			if ((~soc_edid_storage)) begin
				vns_edid_next_state <= 1'd0;
			end
		end
		3'd7: begin
			soc_edid_zero_drv <= 1'd1;
			if (soc_edid_scl_i) begin
				vns_edid_next_state <= 4'd8;
			end
			if (soc_edid_start) begin
				vns_edid_next_state <= 1'd1;
			end
			if ((~soc_edid_storage)) begin
				vns_edid_next_state <= 1'd0;
			end
		end
		4'd8: begin
			soc_edid_zero_drv <= 1'd1;
			if ((~soc_edid_scl_i)) begin
				vns_edid_next_state <= 1'd1;
			end
			if (soc_edid_start) begin
				vns_edid_next_state <= 1'd1;
			end
			if ((~soc_edid_storage)) begin
				vns_edid_next_state <= 1'd0;
			end
		end
		4'd9: begin
			if ((~soc_edid_scl_i)) begin
				if ((soc_edid_counter == 4'd8)) begin
					soc_edid_data_drv_stop <= 1'd1;
					vns_edid_next_state <= 4'd10;
				end else begin
					soc_edid_data_drv_en <= 1'd1;
				end
			end
			if (soc_edid_start) begin
				vns_edid_next_state <= 1'd1;
			end
			if ((~soc_edid_storage)) begin
				vns_edid_next_state <= 1'd0;
			end
		end
		4'd10: begin
			if (soc_edid_scl_rising) begin
				soc_edid_oc_inc <= 1'd1;
				if (soc_edid_sda_i) begin
					vns_edid_next_state <= 1'd0;
				end else begin
					vns_edid_next_state <= 4'd9;
				end
			end
			if (soc_edid_start) begin
				vns_edid_next_state <= 1'd1;
			end
			if ((~soc_edid_storage)) begin
				vns_edid_next_state <= 1'd0;
			end
		end
		default: begin
			if (soc_edid_start) begin
				vns_edid_next_state <= 1'd1;
			end
			if ((~soc_edid_storage)) begin
				vns_edid_next_state <= 1'd0;
			end
		end
	endcase
end
assign soc_locked_status = soc_locked;
assign soc_s7datacapture0_serdes_m_d = soc_s7datacapture0_serdes_m_q;
assign soc_s7datacapture0_serdes_s_d = soc_s7datacapture0_serdes_s_q;
assign soc_s7datacapture0_gearbox_i = soc_s7datacapture0_serdes_m_d;
assign soc_s7datacapture0_d = soc_s7datacapture0_gearbox_o;
assign soc_s7datacapture0_mdata = soc_s7datacapture0_serdes_m_d;
assign soc_s7datacapture0_sdata = (~soc_s7datacapture0_serdes_s_d);
assign soc_s7datacapture0_too_late = (soc_s7datacapture0_lateness == 8'd255);
assign soc_s7datacapture0_too_early = (soc_s7datacapture0_lateness == 1'd0);
assign soc_s7datacapture0_delay_rst = soc_s7datacapture0_do_delay_rst_o;
assign soc_s7datacapture0_delay_master_inc = soc_s7datacapture0_do_delay_master_inc_o;
assign soc_s7datacapture0_delay_master_ce = (soc_s7datacapture0_do_delay_master_inc_o | soc_s7datacapture0_do_delay_master_dec_o);
assign soc_s7datacapture0_delay_slave_inc = soc_s7datacapture0_do_delay_slave_inc_o;
assign soc_s7datacapture0_delay_slave_ce = (soc_s7datacapture0_do_delay_slave_inc_o | soc_s7datacapture0_do_delay_slave_dec_o);
assign soc_s7datacapture0_do_delay_rst_i = (soc_s7datacapture0_dly_ctl_re & soc_s7datacapture0_dly_ctl_r[0]);
assign soc_s7datacapture0_do_delay_master_inc_i = (soc_s7datacapture0_dly_ctl_re & soc_s7datacapture0_dly_ctl_r[1]);
assign soc_s7datacapture0_do_delay_master_dec_i = (soc_s7datacapture0_dly_ctl_re & soc_s7datacapture0_dly_ctl_r[2]);
assign soc_s7datacapture0_do_delay_slave_inc_i = (soc_s7datacapture0_dly_ctl_re & soc_s7datacapture0_dly_ctl_r[3]);
assign soc_s7datacapture0_do_delay_slave_dec_i = (soc_s7datacapture0_dly_ctl_re & soc_s7datacapture0_dly_ctl_r[4]);
assign soc_s7datacapture0_reset_lateness = soc_s7datacapture0_do_reset_lateness_o;
assign soc_s7datacapture0_do_reset_lateness_i = soc_s7datacapture0_phase_reset_re;
assign soc_s7datacapture0_gearbox_rst = (pix1p25x_rst | hdmi_in0_pix_rst);
assign data0_cap_write_clk = pix1p25x_clk;
assign data0_cap_read_clk = hdmi_in0_pix_clk;
assign data0_cap_write_rst = soc_s7datacapture0_gearbox_rst;
assign data0_cap_read_rst = soc_s7datacapture0_gearbox_rst;
assign soc_s7datacapture0_transition = (soc_s7datacapture0_mdata_d != soc_s7datacapture0_mdata);
assign soc_s7datacapture0_inc = (soc_s7datacapture0_transition & (soc_s7datacapture0_mdata == soc_s7datacapture0_sdata));
assign soc_s7datacapture0_dec = (soc_s7datacapture0_transition & (soc_s7datacapture0_mdata != soc_s7datacapture0_sdata));
assign soc_s7datacapture0_do_delay_rst_o = (soc_s7datacapture0_do_delay_rst_toggle_o ^ soc_s7datacapture0_do_delay_rst_toggle_o_r);
assign soc_s7datacapture0_do_delay_master_inc_o = (soc_s7datacapture0_do_delay_master_inc_toggle_o ^ soc_s7datacapture0_do_delay_master_inc_toggle_o_r);
assign soc_s7datacapture0_do_delay_master_dec_o = (soc_s7datacapture0_do_delay_master_dec_toggle_o ^ soc_s7datacapture0_do_delay_master_dec_toggle_o_r);
assign soc_s7datacapture0_do_delay_slave_inc_o = (soc_s7datacapture0_do_delay_slave_inc_toggle_o ^ soc_s7datacapture0_do_delay_slave_inc_toggle_o_r);
assign soc_s7datacapture0_do_delay_slave_dec_o = (soc_s7datacapture0_do_delay_slave_dec_toggle_o ^ soc_s7datacapture0_do_delay_slave_dec_toggle_o_r);
assign soc_s7datacapture0_do_reset_lateness_o = (soc_s7datacapture0_do_reset_lateness_toggle_o ^ soc_s7datacapture0_do_reset_lateness_toggle_o_r);
assign soc_charsync0_raw = {soc_charsync0_raw_data, soc_charsync0_raw_data1};
always @(*) begin
	soc_wer0_transitions <= 8'd0;
	soc_wer0_transitions[0] <= (soc_wer0_data_r[0] ^ soc_wer0_data_r[1]);
	soc_wer0_transitions[1] <= (soc_wer0_data_r[1] ^ soc_wer0_data_r[2]);
	soc_wer0_transitions[2] <= (soc_wer0_data_r[2] ^ soc_wer0_data_r[3]);
	soc_wer0_transitions[3] <= (soc_wer0_data_r[3] ^ soc_wer0_data_r[4]);
	soc_wer0_transitions[4] <= (soc_wer0_data_r[4] ^ soc_wer0_data_r[5]);
	soc_wer0_transitions[5] <= (soc_wer0_data_r[5] ^ soc_wer0_data_r[6]);
	soc_wer0_transitions[6] <= (soc_wer0_data_r[6] ^ soc_wer0_data_r[7]);
	soc_wer0_transitions[7] <= (soc_wer0_data_r[7] ^ soc_wer0_data_r[8]);
end
assign soc_wer0_i = soc_wer0_wer_counter_r_updated;
assign soc_wer0_o = (soc_wer0_toggle_o ^ soc_wer0_toggle_o_r);
assign soc_s7datacapture1_serdes_m_d = soc_s7datacapture1_serdes_m_q;
assign soc_s7datacapture1_serdes_s_d = soc_s7datacapture1_serdes_s_q;
assign soc_s7datacapture1_gearbox_i = soc_s7datacapture1_serdes_m_d;
assign soc_s7datacapture1_d = soc_s7datacapture1_gearbox_o;
assign soc_s7datacapture1_mdata = soc_s7datacapture1_serdes_m_d;
assign soc_s7datacapture1_sdata = (~soc_s7datacapture1_serdes_s_d);
assign soc_s7datacapture1_too_late = (soc_s7datacapture1_lateness == 8'd255);
assign soc_s7datacapture1_too_early = (soc_s7datacapture1_lateness == 1'd0);
assign soc_s7datacapture1_delay_rst = soc_s7datacapture1_do_delay_rst_o;
assign soc_s7datacapture1_delay_master_inc = soc_s7datacapture1_do_delay_master_inc_o;
assign soc_s7datacapture1_delay_master_ce = (soc_s7datacapture1_do_delay_master_inc_o | soc_s7datacapture1_do_delay_master_dec_o);
assign soc_s7datacapture1_delay_slave_inc = soc_s7datacapture1_do_delay_slave_inc_o;
assign soc_s7datacapture1_delay_slave_ce = (soc_s7datacapture1_do_delay_slave_inc_o | soc_s7datacapture1_do_delay_slave_dec_o);
assign soc_s7datacapture1_do_delay_rst_i = (soc_s7datacapture1_dly_ctl_re & soc_s7datacapture1_dly_ctl_r[0]);
assign soc_s7datacapture1_do_delay_master_inc_i = (soc_s7datacapture1_dly_ctl_re & soc_s7datacapture1_dly_ctl_r[1]);
assign soc_s7datacapture1_do_delay_master_dec_i = (soc_s7datacapture1_dly_ctl_re & soc_s7datacapture1_dly_ctl_r[2]);
assign soc_s7datacapture1_do_delay_slave_inc_i = (soc_s7datacapture1_dly_ctl_re & soc_s7datacapture1_dly_ctl_r[3]);
assign soc_s7datacapture1_do_delay_slave_dec_i = (soc_s7datacapture1_dly_ctl_re & soc_s7datacapture1_dly_ctl_r[4]);
assign soc_s7datacapture1_reset_lateness = soc_s7datacapture1_do_reset_lateness_o;
assign soc_s7datacapture1_do_reset_lateness_i = soc_s7datacapture1_phase_reset_re;
assign soc_s7datacapture1_gearbox_rst = (pix1p25x_rst | hdmi_in0_pix_rst);
assign data1_cap_write_clk = pix1p25x_clk;
assign data1_cap_read_clk = hdmi_in0_pix_clk;
assign data1_cap_write_rst = soc_s7datacapture1_gearbox_rst;
assign data1_cap_read_rst = soc_s7datacapture1_gearbox_rst;
assign soc_s7datacapture1_transition = (soc_s7datacapture1_mdata_d != soc_s7datacapture1_mdata);
assign soc_s7datacapture1_inc = (soc_s7datacapture1_transition & (soc_s7datacapture1_mdata == soc_s7datacapture1_sdata));
assign soc_s7datacapture1_dec = (soc_s7datacapture1_transition & (soc_s7datacapture1_mdata != soc_s7datacapture1_sdata));
assign soc_s7datacapture1_do_delay_rst_o = (soc_s7datacapture1_do_delay_rst_toggle_o ^ soc_s7datacapture1_do_delay_rst_toggle_o_r);
assign soc_s7datacapture1_do_delay_master_inc_o = (soc_s7datacapture1_do_delay_master_inc_toggle_o ^ soc_s7datacapture1_do_delay_master_inc_toggle_o_r);
assign soc_s7datacapture1_do_delay_master_dec_o = (soc_s7datacapture1_do_delay_master_dec_toggle_o ^ soc_s7datacapture1_do_delay_master_dec_toggle_o_r);
assign soc_s7datacapture1_do_delay_slave_inc_o = (soc_s7datacapture1_do_delay_slave_inc_toggle_o ^ soc_s7datacapture1_do_delay_slave_inc_toggle_o_r);
assign soc_s7datacapture1_do_delay_slave_dec_o = (soc_s7datacapture1_do_delay_slave_dec_toggle_o ^ soc_s7datacapture1_do_delay_slave_dec_toggle_o_r);
assign soc_s7datacapture1_do_reset_lateness_o = (soc_s7datacapture1_do_reset_lateness_toggle_o ^ soc_s7datacapture1_do_reset_lateness_toggle_o_r);
assign soc_charsync1_raw = {soc_charsync1_raw_data, soc_charsync1_raw_data1};
always @(*) begin
	soc_wer1_transitions <= 8'd0;
	soc_wer1_transitions[0] <= (soc_wer1_data_r[0] ^ soc_wer1_data_r[1]);
	soc_wer1_transitions[1] <= (soc_wer1_data_r[1] ^ soc_wer1_data_r[2]);
	soc_wer1_transitions[2] <= (soc_wer1_data_r[2] ^ soc_wer1_data_r[3]);
	soc_wer1_transitions[3] <= (soc_wer1_data_r[3] ^ soc_wer1_data_r[4]);
	soc_wer1_transitions[4] <= (soc_wer1_data_r[4] ^ soc_wer1_data_r[5]);
	soc_wer1_transitions[5] <= (soc_wer1_data_r[5] ^ soc_wer1_data_r[6]);
	soc_wer1_transitions[6] <= (soc_wer1_data_r[6] ^ soc_wer1_data_r[7]);
	soc_wer1_transitions[7] <= (soc_wer1_data_r[7] ^ soc_wer1_data_r[8]);
end
assign soc_wer1_i = soc_wer1_wer_counter_r_updated;
assign soc_wer1_o = (soc_wer1_toggle_o ^ soc_wer1_toggle_o_r);
assign soc_s7datacapture2_serdes_m_d = soc_s7datacapture2_serdes_m_q;
assign soc_s7datacapture2_serdes_s_d = soc_s7datacapture2_serdes_s_q;
assign soc_s7datacapture2_gearbox_i = soc_s7datacapture2_serdes_m_d;
assign soc_s7datacapture2_d = soc_s7datacapture2_gearbox_o;
assign soc_s7datacapture2_mdata = soc_s7datacapture2_serdes_m_d;
assign soc_s7datacapture2_sdata = (~soc_s7datacapture2_serdes_s_d);
assign soc_s7datacapture2_too_late = (soc_s7datacapture2_lateness == 8'd255);
assign soc_s7datacapture2_too_early = (soc_s7datacapture2_lateness == 1'd0);
assign soc_s7datacapture2_delay_rst = soc_s7datacapture2_do_delay_rst_o;
assign soc_s7datacapture2_delay_master_inc = soc_s7datacapture2_do_delay_master_inc_o;
assign soc_s7datacapture2_delay_master_ce = (soc_s7datacapture2_do_delay_master_inc_o | soc_s7datacapture2_do_delay_master_dec_o);
assign soc_s7datacapture2_delay_slave_inc = soc_s7datacapture2_do_delay_slave_inc_o;
assign soc_s7datacapture2_delay_slave_ce = (soc_s7datacapture2_do_delay_slave_inc_o | soc_s7datacapture2_do_delay_slave_dec_o);
assign soc_s7datacapture2_do_delay_rst_i = (soc_s7datacapture2_dly_ctl_re & soc_s7datacapture2_dly_ctl_r[0]);
assign soc_s7datacapture2_do_delay_master_inc_i = (soc_s7datacapture2_dly_ctl_re & soc_s7datacapture2_dly_ctl_r[1]);
assign soc_s7datacapture2_do_delay_master_dec_i = (soc_s7datacapture2_dly_ctl_re & soc_s7datacapture2_dly_ctl_r[2]);
assign soc_s7datacapture2_do_delay_slave_inc_i = (soc_s7datacapture2_dly_ctl_re & soc_s7datacapture2_dly_ctl_r[3]);
assign soc_s7datacapture2_do_delay_slave_dec_i = (soc_s7datacapture2_dly_ctl_re & soc_s7datacapture2_dly_ctl_r[4]);
assign soc_s7datacapture2_reset_lateness = soc_s7datacapture2_do_reset_lateness_o;
assign soc_s7datacapture2_do_reset_lateness_i = soc_s7datacapture2_phase_reset_re;
assign soc_s7datacapture2_gearbox_rst = (pix1p25x_rst | hdmi_in0_pix_rst);
assign data2_cap_write_clk = pix1p25x_clk;
assign data2_cap_read_clk = hdmi_in0_pix_clk;
assign data2_cap_write_rst = soc_s7datacapture2_gearbox_rst;
assign data2_cap_read_rst = soc_s7datacapture2_gearbox_rst;
assign soc_s7datacapture2_transition = (soc_s7datacapture2_mdata_d != soc_s7datacapture2_mdata);
assign soc_s7datacapture2_inc = (soc_s7datacapture2_transition & (soc_s7datacapture2_mdata == soc_s7datacapture2_sdata));
assign soc_s7datacapture2_dec = (soc_s7datacapture2_transition & (soc_s7datacapture2_mdata != soc_s7datacapture2_sdata));
assign soc_s7datacapture2_do_delay_rst_o = (soc_s7datacapture2_do_delay_rst_toggle_o ^ soc_s7datacapture2_do_delay_rst_toggle_o_r);
assign soc_s7datacapture2_do_delay_master_inc_o = (soc_s7datacapture2_do_delay_master_inc_toggle_o ^ soc_s7datacapture2_do_delay_master_inc_toggle_o_r);
assign soc_s7datacapture2_do_delay_master_dec_o = (soc_s7datacapture2_do_delay_master_dec_toggle_o ^ soc_s7datacapture2_do_delay_master_dec_toggle_o_r);
assign soc_s7datacapture2_do_delay_slave_inc_o = (soc_s7datacapture2_do_delay_slave_inc_toggle_o ^ soc_s7datacapture2_do_delay_slave_inc_toggle_o_r);
assign soc_s7datacapture2_do_delay_slave_dec_o = (soc_s7datacapture2_do_delay_slave_dec_toggle_o ^ soc_s7datacapture2_do_delay_slave_dec_toggle_o_r);
assign soc_s7datacapture2_do_reset_lateness_o = (soc_s7datacapture2_do_reset_lateness_toggle_o ^ soc_s7datacapture2_do_reset_lateness_toggle_o_r);
assign soc_charsync2_raw = {soc_charsync2_raw_data, soc_charsync2_raw_data1};
always @(*) begin
	soc_wer2_transitions <= 8'd0;
	soc_wer2_transitions[0] <= (soc_wer2_data_r[0] ^ soc_wer2_data_r[1]);
	soc_wer2_transitions[1] <= (soc_wer2_data_r[1] ^ soc_wer2_data_r[2]);
	soc_wer2_transitions[2] <= (soc_wer2_data_r[2] ^ soc_wer2_data_r[3]);
	soc_wer2_transitions[3] <= (soc_wer2_data_r[3] ^ soc_wer2_data_r[4]);
	soc_wer2_transitions[4] <= (soc_wer2_data_r[4] ^ soc_wer2_data_r[5]);
	soc_wer2_transitions[5] <= (soc_wer2_data_r[5] ^ soc_wer2_data_r[6]);
	soc_wer2_transitions[6] <= (soc_wer2_data_r[6] ^ soc_wer2_data_r[7]);
	soc_wer2_transitions[7] <= (soc_wer2_data_r[7] ^ soc_wer2_data_r[8]);
end
assign soc_wer2_i = soc_wer2_wer_counter_r_updated;
assign soc_wer2_o = (soc_wer2_toggle_o ^ soc_wer2_toggle_o_r);
assign soc_chansync_syncbuffer0_din = {soc_chansync_data_in0_de, soc_chansync_data_in0_c, soc_chansync_data_in0_d};
assign {soc_chansync_data_out0_de, soc_chansync_data_out0_c, soc_chansync_data_out0_d} = soc_chansync_syncbuffer0_dout;
assign soc_chansync_is_control0 = (~soc_chansync_data_out0_de);
assign soc_chansync_syncbuffer0_re = ((~soc_chansync_is_control0) | soc_chansync_all_control);
assign soc_chansync_syncbuffer1_din = {soc_chansync_data_in1_de, soc_chansync_data_in1_c, soc_chansync_data_in1_d};
assign {soc_chansync_data_out1_de, soc_chansync_data_out1_c, soc_chansync_data_out1_d} = soc_chansync_syncbuffer1_dout;
assign soc_chansync_is_control1 = (~soc_chansync_data_out1_de);
assign soc_chansync_syncbuffer1_re = ((~soc_chansync_is_control1) | soc_chansync_all_control);
assign soc_chansync_syncbuffer2_din = {soc_chansync_data_in2_de, soc_chansync_data_in2_c, soc_chansync_data_in2_d};
assign {soc_chansync_data_out2_de, soc_chansync_data_out2_c, soc_chansync_data_out2_d} = soc_chansync_syncbuffer2_dout;
assign soc_chansync_is_control2 = (~soc_chansync_data_out2_de);
assign soc_chansync_syncbuffer2_re = ((~soc_chansync_is_control2) | soc_chansync_all_control);
assign soc_chansync_all_control = ((soc_chansync_is_control0 & soc_chansync_is_control1) & soc_chansync_is_control2);
assign soc_chansync_some_control = ((soc_chansync_is_control0 | soc_chansync_is_control1) | soc_chansync_is_control2);
assign soc_chansync_syncbuffer0_wrport_adr = soc_chansync_syncbuffer0_produce;
assign soc_chansync_syncbuffer0_wrport_dat_w = soc_chansync_syncbuffer0_din;
assign soc_chansync_syncbuffer0_wrport_we = 1'd1;
assign soc_chansync_syncbuffer0_rdport_adr = soc_chansync_syncbuffer0_consume;
assign soc_chansync_syncbuffer0_dout = soc_chansync_syncbuffer0_rdport_dat_r;
assign soc_chansync_syncbuffer1_wrport_adr = soc_chansync_syncbuffer1_produce;
assign soc_chansync_syncbuffer1_wrport_dat_w = soc_chansync_syncbuffer1_din;
assign soc_chansync_syncbuffer1_wrport_we = 1'd1;
assign soc_chansync_syncbuffer1_rdport_adr = soc_chansync_syncbuffer1_consume;
assign soc_chansync_syncbuffer1_dout = soc_chansync_syncbuffer1_rdport_dat_r;
assign soc_chansync_syncbuffer2_wrport_adr = soc_chansync_syncbuffer2_produce;
assign soc_chansync_syncbuffer2_wrport_dat_w = soc_chansync_syncbuffer2_din;
assign soc_chansync_syncbuffer2_wrport_we = 1'd1;
assign soc_chansync_syncbuffer2_rdport_adr = soc_chansync_syncbuffer2_consume;
assign soc_chansync_syncbuffer2_dout = soc_chansync_syncbuffer2_rdport_dat_r;
assign soc_syncpol_de = soc_syncpol_de_r;
assign soc_syncpol_hsync = soc_syncpol_c_out[0];
assign soc_syncpol_vsync = soc_syncpol_c_out[1];
assign soc_resdetection_pn_de = ((~soc_resdetection_de) & soc_resdetection_de_r);
assign soc_resdetection_p_vsync = (soc_resdetection_vsync & (~soc_resdetection_vsync_r));
assign soc_frame_rgb2ycbcr_sink_valid = soc_frame_valid_i;
assign soc_frame_rgb2ycbcr_sink_payload_r = soc_frame_r;
assign soc_frame_rgb2ycbcr_sink_payload_g = soc_frame_g;
assign soc_frame_rgb2ycbcr_sink_payload_b = soc_frame_b;
assign soc_frame_chroma_downsampler_sink_valid = soc_frame_rgb2ycbcr_source_valid;
assign soc_frame_rgb2ycbcr_source_ready = soc_frame_chroma_downsampler_sink_ready;
assign soc_frame_chroma_downsampler_sink_first = soc_frame_rgb2ycbcr_source_first;
assign soc_frame_chroma_downsampler_sink_last = soc_frame_rgb2ycbcr_source_last;
assign soc_frame_chroma_downsampler_sink_payload_y = soc_frame_rgb2ycbcr_source_payload_y;
assign soc_frame_chroma_downsampler_sink_payload_cb = soc_frame_rgb2ycbcr_source_payload_cb;
assign soc_frame_chroma_downsampler_sink_payload_cr = soc_frame_rgb2ycbcr_source_payload_cr;
assign soc_frame_chroma_downsampler_source_ready = 1'd1;
assign soc_frame_chroma_downsampler_first = (soc_frame_de & (~soc_frame_de_r));
assign soc_frame_new_frame = (soc_frame_next_vsync10 & (~soc_frame_vsync_r));
assign soc_frame_encoded_pixel = {soc_frame_chroma_downsampler_source_payload_cb_cr, soc_frame_chroma_downsampler_source_payload_y};
assign soc_frame_fifo_sink_payload_pixels = soc_frame_cur_word;
assign soc_frame_fifo_sink_valid = soc_frame_cur_word_valid;
assign soc_frame_frame_valid = soc_frame_fifo_source_valid;
assign soc_frame_fifo_source_ready = soc_frame_frame_ready;
assign soc_frame_frame_first = soc_frame_fifo_source_first;
assign soc_frame_frame_last = soc_frame_fifo_source_last;
assign soc_frame_frame_payload_sof = soc_frame_fifo_source_payload_sof;
assign soc_frame_frame_payload_pixels = soc_frame_fifo_source_payload_pixels;
assign soc_frame_busy = 1'd0;
assign soc_frame_pix_overflow_reset = soc_frame_overflow_reset_o;
assign soc_frame_overflow_reset_ack_i = soc_frame_pix_overflow_reset;
assign soc_frame_overflow_w = (soc_frame_sys_overflow & (~soc_frame_overflow_mask));
assign soc_frame_overflow_reset_i = soc_frame_overflow_re;
assign soc_frame_rgb2ycbcr_pipe_ce = (soc_frame_rgb2ycbcr_source_ready | (~soc_frame_rgb2ycbcr_valid_n7));
assign soc_frame_rgb2ycbcr_sink_ready = soc_frame_rgb2ycbcr_pipe_ce;
assign soc_frame_rgb2ycbcr_source_valid = soc_frame_rgb2ycbcr_valid_n7;
assign soc_frame_rgb2ycbcr_busy = ((((((((1'd0 | soc_frame_rgb2ycbcr_valid_n0) | soc_frame_rgb2ycbcr_valid_n1) | soc_frame_rgb2ycbcr_valid_n2) | soc_frame_rgb2ycbcr_valid_n3) | soc_frame_rgb2ycbcr_valid_n4) | soc_frame_rgb2ycbcr_valid_n5) | soc_frame_rgb2ycbcr_valid_n6) | soc_frame_rgb2ycbcr_valid_n7);
assign soc_frame_rgb2ycbcr_source_first = soc_frame_rgb2ycbcr_first_n7;
assign soc_frame_rgb2ycbcr_source_last = soc_frame_rgb2ycbcr_last_n7;
assign soc_frame_rgb2ycbcr_ce = soc_frame_rgb2ycbcr_pipe_ce;
assign soc_frame_rgb2ycbcr_sink_r = soc_frame_rgb2ycbcr_sink_payload_r;
assign soc_frame_rgb2ycbcr_sink_g = soc_frame_rgb2ycbcr_sink_payload_g;
assign soc_frame_rgb2ycbcr_sink_b = soc_frame_rgb2ycbcr_sink_payload_b;
assign soc_frame_rgb2ycbcr_source_payload_y = soc_frame_rgb2ycbcr_source_y;
assign soc_frame_rgb2ycbcr_source_payload_cb = soc_frame_rgb2ycbcr_source_cb;
assign soc_frame_rgb2ycbcr_source_payload_cr = soc_frame_rgb2ycbcr_source_cr;
assign soc_frame_chroma_downsampler_pipe_ce = (soc_frame_chroma_downsampler_source_ready | (~soc_frame_chroma_downsampler_valid_n2));
assign soc_frame_chroma_downsampler_sink_ready = soc_frame_chroma_downsampler_pipe_ce;
assign soc_frame_chroma_downsampler_source_valid = soc_frame_chroma_downsampler_valid_n2;
assign soc_frame_chroma_downsampler_busy = (((1'd0 | soc_frame_chroma_downsampler_valid_n0) | soc_frame_chroma_downsampler_valid_n1) | soc_frame_chroma_downsampler_valid_n2);
assign soc_frame_chroma_downsampler_source_first = soc_frame_chroma_downsampler_first_n2;
assign soc_frame_chroma_downsampler_source_last = soc_frame_chroma_downsampler_last_n2;
assign soc_frame_chroma_downsampler_ce = soc_frame_chroma_downsampler_pipe_ce;
assign soc_frame_chroma_downsampler_sink_y = soc_frame_chroma_downsampler_sink_payload_y;
assign soc_frame_chroma_downsampler_sink_cb = soc_frame_chroma_downsampler_sink_payload_cb;
assign soc_frame_chroma_downsampler_sink_cr = soc_frame_chroma_downsampler_sink_payload_cr;
assign soc_frame_chroma_downsampler_source_payload_y = soc_frame_chroma_downsampler_source_y;
assign soc_frame_chroma_downsampler_source_payload_cb_cr = soc_frame_chroma_downsampler_source_cb_cr;
assign soc_frame_chroma_downsampler_cb_mean = soc_frame_chroma_downsampler_cb_sum[8:1];
assign soc_frame_chroma_downsampler_cr_mean = soc_frame_chroma_downsampler_cr_sum[8:1];
assign soc_frame_fifo_asyncfifo_din = {soc_frame_fifo_fifo_in_last, soc_frame_fifo_fifo_in_first, soc_frame_fifo_fifo_in_payload_pixels, soc_frame_fifo_fifo_in_payload_sof};
assign {soc_frame_fifo_fifo_out_last, soc_frame_fifo_fifo_out_first, soc_frame_fifo_fifo_out_payload_pixels, soc_frame_fifo_fifo_out_payload_sof} = soc_frame_fifo_asyncfifo_dout;
assign soc_frame_fifo_sink_ready = soc_frame_fifo_asyncfifo_writable;
assign soc_frame_fifo_asyncfifo_we = soc_frame_fifo_sink_valid;
assign soc_frame_fifo_fifo_in_first = soc_frame_fifo_sink_first;
assign soc_frame_fifo_fifo_in_last = soc_frame_fifo_sink_last;
assign soc_frame_fifo_fifo_in_payload_sof = soc_frame_fifo_sink_payload_sof;
assign soc_frame_fifo_fifo_in_payload_pixels = soc_frame_fifo_sink_payload_pixels;
assign soc_frame_fifo_source_valid = soc_frame_fifo_asyncfifo_readable;
assign soc_frame_fifo_source_first = soc_frame_fifo_fifo_out_first;
assign soc_frame_fifo_source_last = soc_frame_fifo_fifo_out_last;
assign soc_frame_fifo_source_payload_sof = soc_frame_fifo_fifo_out_payload_sof;
assign soc_frame_fifo_source_payload_pixels = soc_frame_fifo_fifo_out_payload_pixels;
assign soc_frame_fifo_asyncfifo_re = soc_frame_fifo_source_ready;
assign soc_frame_fifo_graycounter0_ce = (soc_frame_fifo_asyncfifo_writable & soc_frame_fifo_asyncfifo_we);
assign soc_frame_fifo_graycounter1_ce = (soc_frame_fifo_asyncfifo_readable & soc_frame_fifo_asyncfifo_re);
assign soc_frame_fifo_asyncfifo_writable = (((soc_frame_fifo_graycounter0_q[9] == soc_frame_fifo_consume_wdomain[9]) | (soc_frame_fifo_graycounter0_q[8] == soc_frame_fifo_consume_wdomain[8])) | (soc_frame_fifo_graycounter0_q[7:0] != soc_frame_fifo_consume_wdomain[7:0]));
assign soc_frame_fifo_asyncfifo_readable = (soc_frame_fifo_graycounter1_q != soc_frame_fifo_produce_rdomain);
assign soc_frame_fifo_wrport_adr = soc_frame_fifo_graycounter0_q_binary[8:0];
assign soc_frame_fifo_wrport_dat_w = soc_frame_fifo_asyncfifo_din;
assign soc_frame_fifo_wrport_we = soc_frame_fifo_graycounter0_ce;
assign soc_frame_fifo_rdport_adr = soc_frame_fifo_graycounter1_q_next_binary[8:0];
assign soc_frame_fifo_asyncfifo_dout = soc_frame_fifo_rdport_dat_r;
always @(*) begin
	soc_frame_fifo_graycounter0_q_next_binary <= 10'd0;
	if (soc_frame_fifo_graycounter0_ce) begin
		soc_frame_fifo_graycounter0_q_next_binary <= (soc_frame_fifo_graycounter0_q_binary + 1'd1);
	end else begin
		soc_frame_fifo_graycounter0_q_next_binary <= soc_frame_fifo_graycounter0_q_binary;
	end
end
assign soc_frame_fifo_graycounter0_q_next = (soc_frame_fifo_graycounter0_q_next_binary ^ soc_frame_fifo_graycounter0_q_next_binary[9:1]);
always @(*) begin
	soc_frame_fifo_graycounter1_q_next_binary <= 10'd0;
	if (soc_frame_fifo_graycounter1_ce) begin
		soc_frame_fifo_graycounter1_q_next_binary <= (soc_frame_fifo_graycounter1_q_binary + 1'd1);
	end else begin
		soc_frame_fifo_graycounter1_q_next_binary <= soc_frame_fifo_graycounter1_q_binary;
	end
end
assign soc_frame_fifo_graycounter1_q_next = (soc_frame_fifo_graycounter1_q_next_binary ^ soc_frame_fifo_graycounter1_q_next_binary[9:1]);
assign soc_frame_overflow_reset_o = (soc_frame_overflow_reset_toggle_o ^ soc_frame_overflow_reset_toggle_o_r);
assign soc_frame_overflow_reset_ack_o = (soc_frame_overflow_reset_ack_toggle_o ^ soc_frame_overflow_reset_ack_toggle_o_r);
assign soc_dma_slot_array_address_reached = soc_dma_current_address;
assign soc_dma_last_word = (soc_dma_mwords_remaining == 1'd1);
assign soc_dma_memory_word = {soc_dma_frame_payload_pixels, soc_dma_frame_payload_pixels, soc_dma_frame_payload_pixels, soc_dma_frame_payload_pixels, soc_dma_frame_payload_pixels, soc_dma_frame_payload_pixels, soc_dma_frame_payload_pixels, soc_dma_frame_payload_pixels};
assign soc_dma_sink_sink_payload_address = soc_dma_current_address;
assign soc_dma_sink_sink_payload_data = soc_dma_memory_word;
assign soc_dma_slot_array_change_slot = ((~soc_dma_slot_array_address_valid) | soc_dma_slot_array_address_done);
assign soc_dma_slot_array_address = vns_comb_rhs_array_muxed36;
assign soc_dma_slot_array_address_valid = vns_comb_rhs_array_muxed37;
assign soc_dma_slot_array_slot0_address_reached = soc_dma_slot_array_address_reached;
assign soc_dma_slot_array_slot1_address_reached = soc_dma_slot_array_address_reached;
assign soc_dma_slot_array_slot0_address_done = (soc_dma_slot_array_address_done & (soc_dma_slot_array_current_slot == 1'd0));
assign soc_dma_slot_array_slot1_address_done = (soc_dma_slot_array_address_done & (soc_dma_slot_array_current_slot == 1'd1));
always @(*) begin
	soc_dma_slot_array_slot0_clear <= 1'd0;
	if ((soc_dma_slot_array_pending_re & soc_dma_slot_array_pending_r[0])) begin
		soc_dma_slot_array_slot0_clear <= 1'd1;
	end
end
always @(*) begin
	soc_dma_slot_array_status_w <= 2'd0;
	soc_dma_slot_array_status_w[0] <= soc_dma_slot_array_slot0_status;
	soc_dma_slot_array_status_w[1] <= soc_dma_slot_array_slot1_status;
end
always @(*) begin
	soc_dma_slot_array_slot1_clear <= 1'd0;
	if ((soc_dma_slot_array_pending_re & soc_dma_slot_array_pending_r[1])) begin
		soc_dma_slot_array_slot1_clear <= 1'd1;
	end
end
always @(*) begin
	soc_dma_slot_array_pending_w <= 2'd0;
	soc_dma_slot_array_pending_w[0] <= soc_dma_slot_array_slot0_pending;
	soc_dma_slot_array_pending_w[1] <= soc_dma_slot_array_slot1_pending;
end
assign soc_dma_slot_array_irq = ((soc_dma_slot_array_pending_w[0] & soc_dma_slot_array_storage[0]) | (soc_dma_slot_array_pending_w[1] & soc_dma_slot_array_storage[1]));
assign soc_dma_slot_array_slot0_status = soc_dma_slot_array_slot0_trigger;
assign soc_dma_slot_array_slot0_pending = soc_dma_slot_array_slot0_trigger;
assign soc_dma_slot_array_slot1_status = soc_dma_slot_array_slot1_trigger;
assign soc_dma_slot_array_slot1_pending = soc_dma_slot_array_slot1_trigger;
assign soc_dma_slot_array_slot0_address = soc_dma_slot_array_slot0_address_storage;
assign soc_dma_slot_array_slot0_address_valid = soc_dma_slot_array_slot0_status_storage[0];
assign soc_dma_slot_array_slot0_status_dat_w = 2'd2;
assign soc_dma_slot_array_slot0_status_we = soc_dma_slot_array_slot0_address_done;
assign soc_dma_slot_array_slot0_address_dat_w = soc_dma_slot_array_slot0_address_reached;
assign soc_dma_slot_array_slot0_address_we = soc_dma_slot_array_slot0_address_done;
assign soc_dma_slot_array_slot0_trigger = soc_dma_slot_array_slot0_status_storage[1];
assign soc_dma_slot_array_slot1_address = soc_dma_slot_array_slot1_address_storage;
assign soc_dma_slot_array_slot1_address_valid = soc_dma_slot_array_slot1_status_storage[0];
assign soc_dma_slot_array_slot1_status_dat_w = 2'd2;
assign soc_dma_slot_array_slot1_status_we = soc_dma_slot_array_slot1_address_done;
assign soc_dma_slot_array_slot1_address_dat_w = soc_dma_slot_array_slot1_address_reached;
assign soc_dma_slot_array_slot1_address_we = soc_dma_slot_array_slot1_address_done;
assign soc_dma_slot_array_slot1_trigger = soc_dma_slot_array_slot1_status_storage[1];
assign soc_litedramcrossbar_cmd_payload_we = 1'd1;
assign soc_litedramcrossbar_cmd_valid = (soc_dma_fifo_sink_ready & soc_dma_sink_sink_valid);
assign soc_litedramcrossbar_cmd_payload_adr = soc_dma_sink_sink_payload_address;
assign soc_dma_sink_sink_ready = (soc_dma_fifo_sink_ready & soc_litedramcrossbar_cmd_ready);
assign soc_dma_fifo_sink_valid = (soc_dma_sink_sink_valid & soc_litedramcrossbar_cmd_ready);
assign soc_dma_fifo_sink_payload_data = soc_dma_sink_sink_payload_data;
assign soc_litedramcrossbar_wdata_valid = soc_dma_fifo_source_valid;
assign soc_dma_fifo_source_ready = soc_litedramcrossbar_wdata_ready;
assign soc_litedramcrossbar_wdata_payload_we = 16'd65535;
assign soc_litedramcrossbar_wdata_payload_data = soc_dma_fifo_source_payload_data;
assign soc_dma_fifo_syncfifo_din = {soc_dma_fifo_fifo_in_last, soc_dma_fifo_fifo_in_first, soc_dma_fifo_fifo_in_payload_data};
assign {soc_dma_fifo_fifo_out_last, soc_dma_fifo_fifo_out_first, soc_dma_fifo_fifo_out_payload_data} = soc_dma_fifo_syncfifo_dout;
assign soc_dma_fifo_sink_ready = soc_dma_fifo_syncfifo_writable;
assign soc_dma_fifo_syncfifo_we = soc_dma_fifo_sink_valid;
assign soc_dma_fifo_fifo_in_first = soc_dma_fifo_sink_first;
assign soc_dma_fifo_fifo_in_last = soc_dma_fifo_sink_last;
assign soc_dma_fifo_fifo_in_payload_data = soc_dma_fifo_sink_payload_data;
assign soc_dma_fifo_source_valid = soc_dma_fifo_syncfifo_readable;
assign soc_dma_fifo_source_first = soc_dma_fifo_fifo_out_first;
assign soc_dma_fifo_source_last = soc_dma_fifo_fifo_out_last;
assign soc_dma_fifo_source_payload_data = soc_dma_fifo_fifo_out_payload_data;
assign soc_dma_fifo_syncfifo_re = soc_dma_fifo_source_ready;
always @(*) begin
	soc_dma_fifo_wrport_adr <= 4'd0;
	if (soc_dma_fifo_replace) begin
		soc_dma_fifo_wrport_adr <= (soc_dma_fifo_produce - 1'd1);
	end else begin
		soc_dma_fifo_wrport_adr <= soc_dma_fifo_produce;
	end
end
assign soc_dma_fifo_wrport_dat_w = soc_dma_fifo_syncfifo_din;
assign soc_dma_fifo_wrport_we = (soc_dma_fifo_syncfifo_we & (soc_dma_fifo_syncfifo_writable | soc_dma_fifo_replace));
assign soc_dma_fifo_do_read = (soc_dma_fifo_syncfifo_readable & soc_dma_fifo_syncfifo_re);
assign soc_dma_fifo_rdport_adr = soc_dma_fifo_consume;
assign soc_dma_fifo_syncfifo_dout = soc_dma_fifo_rdport_dat_r;
assign soc_dma_fifo_syncfifo_writable = (soc_dma_fifo_level != 5'd16);
assign soc_dma_fifo_syncfifo_readable = (soc_dma_fifo_level != 1'd0);
always @(*) begin
	soc_dma_sink_sink_valid <= 1'd0;
	soc_dma_slot_array_address_done <= 1'd0;
	vns_dma_next_state <= 2'd0;
	soc_dma_frame_ready <= 1'd0;
	soc_dma_reset_words <= 1'd0;
	soc_dma_count_word <= 1'd0;
	vns_dma_next_state <= vns_dma_state;
	case (vns_dma_state)
		1'd1: begin
			soc_dma_frame_ready <= soc_dma_sink_sink_ready;
			if (soc_dma_frame_valid) begin
				soc_dma_sink_sink_valid <= 1'd1;
				if (soc_dma_sink_sink_ready) begin
					soc_dma_count_word <= 1'd1;
					if (soc_dma_last_word) begin
						vns_dma_next_state <= 2'd2;
					end
				end
			end
		end
		2'd2: begin
			if ((~soc_litedramcrossbar_wdata_valid)) begin
				soc_dma_slot_array_address_done <= 1'd1;
				vns_dma_next_state <= 1'd0;
			end
		end
		default: begin
			soc_dma_reset_words <= 1'd1;
			soc_dma_frame_ready <= ((~soc_dma_slot_array_address_valid) | (~soc_dma_frame_payload_sof));
			if (((soc_dma_slot_array_address_valid & soc_dma_frame_payload_sof) & soc_dma_frame_valid)) begin
				vns_dma_next_state <= 1'd1;
			end
		end
	endcase
end
assign fmeter_clk = soc_hdmi_in0_freq_clk0;
assign soc_hdmi_in0_freq_period_done = (soc_hdmi_in0_freq_period_counter == 27'd100000000);
assign soc_hdmi_in0_freq_ce = 1'd1;
assign soc_hdmi_in0_freq_sampler_latch = soc_hdmi_in0_freq_period_done;
assign soc_hdmi_in0_freq_sampler_i = soc_hdmi_in0_freq_gray_decoder_o;
assign soc_hdmi_in0_freq_status = soc_hdmi_in0_freq_sampler_o;
always @(*) begin
	soc_hdmi_in0_freq_q_next_binary <= 6'd0;
	if (soc_hdmi_in0_freq_ce) begin
		soc_hdmi_in0_freq_q_next_binary <= (soc_hdmi_in0_freq_q_binary + 1'd1);
	end else begin
		soc_hdmi_in0_freq_q_next_binary <= soc_hdmi_in0_freq_q_binary;
	end
end
assign soc_hdmi_in0_freq_q_next = (soc_hdmi_in0_freq_q_next_binary ^ soc_hdmi_in0_freq_q_next_binary[5:1]);
always @(*) begin
	soc_hdmi_in0_freq_gray_decoder_o_comb <= 6'd0;
	soc_hdmi_in0_freq_gray_decoder_o_comb[5] <= soc_hdmi_in0_freq_gray_decoder_i[5];
	soc_hdmi_in0_freq_gray_decoder_o_comb[4] <= (soc_hdmi_in0_freq_gray_decoder_o_comb[5] ^ soc_hdmi_in0_freq_gray_decoder_i[4]);
	soc_hdmi_in0_freq_gray_decoder_o_comb[3] <= (soc_hdmi_in0_freq_gray_decoder_o_comb[4] ^ soc_hdmi_in0_freq_gray_decoder_i[3]);
	soc_hdmi_in0_freq_gray_decoder_o_comb[2] <= (soc_hdmi_in0_freq_gray_decoder_o_comb[3] ^ soc_hdmi_in0_freq_gray_decoder_i[2]);
	soc_hdmi_in0_freq_gray_decoder_o_comb[1] <= (soc_hdmi_in0_freq_gray_decoder_o_comb[2] ^ soc_hdmi_in0_freq_gray_decoder_i[1]);
	soc_hdmi_in0_freq_gray_decoder_o_comb[0] <= (soc_hdmi_in0_freq_gray_decoder_o_comb[1] ^ soc_hdmi_in0_freq_gray_decoder_i[0]);
end
assign soc_hdmi_in0_freq_sampler_inc = (soc_hdmi_in0_freq_sampler_i - soc_hdmi_in0_freq_sampler_i_d);
assign soc_hdmi_out0_core_source_source_ready = 1'd1;
assign soc_hdmi_out0_resetinserter_reset = (soc_hdmi_out0_core_source_source_param_de & (~soc_hdmi_out0_de_r));
assign soc_hdmi_out0_resetinserter_sink_sink_valid = soc_hdmi_out0_core_source_valid_d;
assign soc_hdmi_out0_resetinserter_sink_sink_payload_y = soc_hdmi_out0_core_source_data_d[7:0];
assign soc_hdmi_out0_resetinserter_sink_sink_payload_cb_cr = soc_hdmi_out0_core_source_data_d[15:8];
assign soc_hdmi_out0_sink_valid = soc_hdmi_out0_resetinserter_source_source_valid;
assign soc_hdmi_out0_resetinserter_source_source_ready = soc_hdmi_out0_sink_ready;
assign soc_hdmi_out0_sink_first = soc_hdmi_out0_resetinserter_source_source_first;
assign soc_hdmi_out0_sink_last = soc_hdmi_out0_resetinserter_source_source_last;
assign soc_hdmi_out0_sink_payload_y = soc_hdmi_out0_resetinserter_source_source_payload_y;
assign soc_hdmi_out0_sink_payload_cb = soc_hdmi_out0_resetinserter_source_source_payload_cb;
assign soc_hdmi_out0_sink_payload_cr = soc_hdmi_out0_resetinserter_source_source_payload_cr;
assign soc_hdmi_out0_driver_sink_sink_valid = soc_hdmi_out0_source_valid;
assign soc_hdmi_out0_source_ready = soc_hdmi_out0_driver_sink_sink_ready;
assign soc_hdmi_out0_driver_sink_sink_first = soc_hdmi_out0_source_first;
assign soc_hdmi_out0_driver_sink_sink_last = soc_hdmi_out0_source_last;
assign soc_hdmi_out0_driver_sink_sink_payload_r = soc_hdmi_out0_source_payload_r;
assign soc_hdmi_out0_driver_sink_sink_payload_g = soc_hdmi_out0_source_payload_g;
assign soc_hdmi_out0_driver_sink_sink_payload_b = soc_hdmi_out0_source_payload_b;
assign soc_hdmi_out0_sink_payload_de = soc_hdmi_out0_core_source_source_param_de;
assign soc_hdmi_out0_sink_payload_vsync = soc_hdmi_out0_core_source_source_param_vsync;
assign soc_hdmi_out0_sink_payload_hsync = soc_hdmi_out0_core_source_source_param_hsync;
assign soc_hdmi_out0_driver_sink_sink_param_de = soc_hdmi_out0_source_payload_de;
assign soc_hdmi_out0_driver_sink_sink_param_vsync = soc_hdmi_out0_source_payload_vsync;
assign soc_hdmi_out0_driver_sink_sink_param_hsync = soc_hdmi_out0_source_payload_hsync;
assign soc_hdmi_out0_core_timinggenerator_sink_valid = soc_hdmi_out0_core_initiator_source_source_valid;
assign soc_hdmi_out0_core_dmareader_sink_valid = soc_hdmi_out0_core_initiator_source_source_valid;
assign soc_hdmi_out0_core_initiator_source_source_ready = soc_hdmi_out0_core_timinggenerator_sink_ready;
assign soc_hdmi_out0_core_source_source_valid = (soc_hdmi_out0_core_timinggenerator_source_valid & ((~soc_hdmi_out0_core_timinggenerator_source_payload_de) | soc_hdmi_out0_core_dmareader_source_valid));
always @(*) begin
	soc_hdmi_out0_core_timinggenerator_source_ready <= 1'd0;
	soc_hdmi_out0_core_dmareader_source_ready <= 1'd0;
	if ((~soc_hdmi_out0_core_initiator_source_source_valid)) begin
		soc_hdmi_out0_core_timinggenerator_source_ready <= 1'd1;
		soc_hdmi_out0_core_dmareader_source_ready <= 1'd1;
	end else begin
		if ((soc_hdmi_out0_core_source_source_valid & soc_hdmi_out0_core_source_source_ready)) begin
			soc_hdmi_out0_core_timinggenerator_source_ready <= 1'd1;
			soc_hdmi_out0_core_dmareader_source_ready <= soc_hdmi_out0_core_timinggenerator_source_payload_de;
		end
	end
end
assign soc_hdmi_out0_core_timinggenerator_sink_payload_hres = soc_hdmi_out0_core_initiator_source_source_payload_hres;
assign soc_hdmi_out0_core_timinggenerator_sink_payload_hsync_start = soc_hdmi_out0_core_initiator_source_source_payload_hsync_start;
assign soc_hdmi_out0_core_timinggenerator_sink_payload_hsync_end = soc_hdmi_out0_core_initiator_source_source_payload_hsync_end;
assign soc_hdmi_out0_core_timinggenerator_sink_payload_hscan = soc_hdmi_out0_core_initiator_source_source_payload_hscan;
assign soc_hdmi_out0_core_timinggenerator_sink_payload_vres = soc_hdmi_out0_core_initiator_source_source_payload_vres;
assign soc_hdmi_out0_core_timinggenerator_sink_payload_vsync_start = soc_hdmi_out0_core_initiator_source_source_payload_vsync_start;
assign soc_hdmi_out0_core_timinggenerator_sink_payload_vsync_end = soc_hdmi_out0_core_initiator_source_source_payload_vsync_end;
assign soc_hdmi_out0_core_timinggenerator_sink_payload_vscan = soc_hdmi_out0_core_initiator_source_source_payload_vscan;
assign soc_hdmi_out0_core_dmareader_sink_payload_base = soc_hdmi_out0_core_initiator_source_source_payload_base;
assign soc_hdmi_out0_core_dmareader_sink_payload_length = soc_hdmi_out0_core_initiator_source_source_payload_length;
assign soc_hdmi_out0_core_source_source_param_de = soc_hdmi_out0_core_timinggenerator_source_payload_de;
assign soc_hdmi_out0_core_source_source_param_hsync = soc_hdmi_out0_core_timinggenerator_source_payload_hsync;
assign soc_hdmi_out0_core_source_source_param_vsync = soc_hdmi_out0_core_timinggenerator_source_payload_vsync;
assign soc_hdmi_out0_core_source_source_payload_data = soc_hdmi_out0_core_dmareader_source_payload_data;
assign soc_hdmi_out0_core_i = soc_hdmi_out0_core_underflow_update_underflow_update_re;
assign soc_hdmi_out0_core_underflow_update = soc_hdmi_out0_core_o;
assign soc_hdmi_out0_core_initiator_cdc_sink_payload_hres = soc_hdmi_out0_core_initiator_csrstorage0_storage;
assign soc_hdmi_out0_core_initiator_cdc_sink_payload_hsync_start = soc_hdmi_out0_core_initiator_csrstorage1_storage;
assign soc_hdmi_out0_core_initiator_cdc_sink_payload_hsync_end = soc_hdmi_out0_core_initiator_csrstorage2_storage;
assign soc_hdmi_out0_core_initiator_cdc_sink_payload_hscan = soc_hdmi_out0_core_initiator_csrstorage3_storage;
assign soc_hdmi_out0_core_initiator_cdc_sink_payload_vres = soc_hdmi_out0_core_initiator_csrstorage4_storage;
assign soc_hdmi_out0_core_initiator_cdc_sink_payload_vsync_start = soc_hdmi_out0_core_initiator_csrstorage5_storage;
assign soc_hdmi_out0_core_initiator_cdc_sink_payload_vsync_end = soc_hdmi_out0_core_initiator_csrstorage6_storage;
assign soc_hdmi_out0_core_initiator_cdc_sink_payload_vscan = soc_hdmi_out0_core_initiator_csrstorage7_storage;
assign soc_hdmi_out0_core_initiator_cdc_sink_payload_base = soc_hdmi_out0_core_initiator_csrstorage8_storage;
assign soc_hdmi_out0_core_initiator_cdc_sink_payload_length = soc_hdmi_out0_core_initiator_csrstorage9_storage;
assign soc_hdmi_out0_core_initiator_cdc_sink_valid = soc_hdmi_out0_core_initiator_enable_storage;
assign soc_hdmi_out0_core_initiator_source_source_valid = soc_hdmi_out0_core_initiator_cdc_source_valid;
assign soc_hdmi_out0_core_initiator_cdc_source_ready = soc_hdmi_out0_core_initiator_source_source_ready;
assign soc_hdmi_out0_core_initiator_source_source_first = soc_hdmi_out0_core_initiator_cdc_source_first;
assign soc_hdmi_out0_core_initiator_source_source_last = soc_hdmi_out0_core_initiator_cdc_source_last;
assign soc_hdmi_out0_core_initiator_source_source_payload_hres = soc_hdmi_out0_core_initiator_cdc_source_payload_hres;
assign soc_hdmi_out0_core_initiator_source_source_payload_hsync_start = soc_hdmi_out0_core_initiator_cdc_source_payload_hsync_start;
assign soc_hdmi_out0_core_initiator_source_source_payload_hsync_end = soc_hdmi_out0_core_initiator_cdc_source_payload_hsync_end;
assign soc_hdmi_out0_core_initiator_source_source_payload_hscan = soc_hdmi_out0_core_initiator_cdc_source_payload_hscan;
assign soc_hdmi_out0_core_initiator_source_source_payload_vres = soc_hdmi_out0_core_initiator_cdc_source_payload_vres;
assign soc_hdmi_out0_core_initiator_source_source_payload_vsync_start = soc_hdmi_out0_core_initiator_cdc_source_payload_vsync_start;
assign soc_hdmi_out0_core_initiator_source_source_payload_vsync_end = soc_hdmi_out0_core_initiator_cdc_source_payload_vsync_end;
assign soc_hdmi_out0_core_initiator_source_source_payload_vscan = soc_hdmi_out0_core_initiator_cdc_source_payload_vscan;
assign soc_hdmi_out0_core_initiator_source_source_payload_base = soc_hdmi_out0_core_initiator_cdc_source_payload_base;
assign soc_hdmi_out0_core_initiator_source_source_payload_length = soc_hdmi_out0_core_initiator_cdc_source_payload_length;
assign soc_hdmi_out0_core_initiator_cdc_asyncfifo_din = {soc_hdmi_out0_core_initiator_cdc_fifo_in_last, soc_hdmi_out0_core_initiator_cdc_fifo_in_first, soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_length, soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_base, soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vscan, soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_end, soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_start, soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vres, soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hscan, soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_end, soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_start, soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hres};
assign {soc_hdmi_out0_core_initiator_cdc_fifo_out_last, soc_hdmi_out0_core_initiator_cdc_fifo_out_first, soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_length, soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_base, soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vscan, soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_end, soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_start, soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vres, soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hscan, soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_end, soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_start, soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hres} = soc_hdmi_out0_core_initiator_cdc_asyncfifo_dout;
assign soc_hdmi_out0_core_initiator_cdc_sink_ready = soc_hdmi_out0_core_initiator_cdc_asyncfifo_writable;
assign soc_hdmi_out0_core_initiator_cdc_asyncfifo_we = soc_hdmi_out0_core_initiator_cdc_sink_valid;
assign soc_hdmi_out0_core_initiator_cdc_fifo_in_first = soc_hdmi_out0_core_initiator_cdc_sink_first;
assign soc_hdmi_out0_core_initiator_cdc_fifo_in_last = soc_hdmi_out0_core_initiator_cdc_sink_last;
assign soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hres = soc_hdmi_out0_core_initiator_cdc_sink_payload_hres;
assign soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_start = soc_hdmi_out0_core_initiator_cdc_sink_payload_hsync_start;
assign soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hsync_end = soc_hdmi_out0_core_initiator_cdc_sink_payload_hsync_end;
assign soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_hscan = soc_hdmi_out0_core_initiator_cdc_sink_payload_hscan;
assign soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vres = soc_hdmi_out0_core_initiator_cdc_sink_payload_vres;
assign soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_start = soc_hdmi_out0_core_initiator_cdc_sink_payload_vsync_start;
assign soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vsync_end = soc_hdmi_out0_core_initiator_cdc_sink_payload_vsync_end;
assign soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_vscan = soc_hdmi_out0_core_initiator_cdc_sink_payload_vscan;
assign soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_base = soc_hdmi_out0_core_initiator_cdc_sink_payload_base;
assign soc_hdmi_out0_core_initiator_cdc_fifo_in_payload_length = soc_hdmi_out0_core_initiator_cdc_sink_payload_length;
assign soc_hdmi_out0_core_initiator_cdc_source_valid = soc_hdmi_out0_core_initiator_cdc_asyncfifo_readable;
assign soc_hdmi_out0_core_initiator_cdc_source_first = soc_hdmi_out0_core_initiator_cdc_fifo_out_first;
assign soc_hdmi_out0_core_initiator_cdc_source_last = soc_hdmi_out0_core_initiator_cdc_fifo_out_last;
assign soc_hdmi_out0_core_initiator_cdc_source_payload_hres = soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hres;
assign soc_hdmi_out0_core_initiator_cdc_source_payload_hsync_start = soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_start;
assign soc_hdmi_out0_core_initiator_cdc_source_payload_hsync_end = soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hsync_end;
assign soc_hdmi_out0_core_initiator_cdc_source_payload_hscan = soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_hscan;
assign soc_hdmi_out0_core_initiator_cdc_source_payload_vres = soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vres;
assign soc_hdmi_out0_core_initiator_cdc_source_payload_vsync_start = soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_start;
assign soc_hdmi_out0_core_initiator_cdc_source_payload_vsync_end = soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vsync_end;
assign soc_hdmi_out0_core_initiator_cdc_source_payload_vscan = soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_vscan;
assign soc_hdmi_out0_core_initiator_cdc_source_payload_base = soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_base;
assign soc_hdmi_out0_core_initiator_cdc_source_payload_length = soc_hdmi_out0_core_initiator_cdc_fifo_out_payload_length;
assign soc_hdmi_out0_core_initiator_cdc_asyncfifo_re = soc_hdmi_out0_core_initiator_cdc_source_ready;
assign soc_hdmi_out0_core_initiator_cdc_graycounter0_ce = (soc_hdmi_out0_core_initiator_cdc_asyncfifo_writable & soc_hdmi_out0_core_initiator_cdc_asyncfifo_we);
assign soc_hdmi_out0_core_initiator_cdc_graycounter1_ce = (soc_hdmi_out0_core_initiator_cdc_asyncfifo_readable & soc_hdmi_out0_core_initiator_cdc_asyncfifo_re);
assign soc_hdmi_out0_core_initiator_cdc_asyncfifo_writable = ((soc_hdmi_out0_core_initiator_cdc_graycounter0_q[1] == soc_hdmi_out0_core_initiator_cdc_consume_wdomain[1]) | (soc_hdmi_out0_core_initiator_cdc_graycounter0_q[0] == soc_hdmi_out0_core_initiator_cdc_consume_wdomain[0]));
assign soc_hdmi_out0_core_initiator_cdc_asyncfifo_readable = (soc_hdmi_out0_core_initiator_cdc_graycounter1_q != soc_hdmi_out0_core_initiator_cdc_produce_rdomain);
assign soc_hdmi_out0_core_initiator_cdc_wrport_adr = soc_hdmi_out0_core_initiator_cdc_graycounter0_q_binary[0];
assign soc_hdmi_out0_core_initiator_cdc_wrport_dat_w = soc_hdmi_out0_core_initiator_cdc_asyncfifo_din;
assign soc_hdmi_out0_core_initiator_cdc_wrport_we = soc_hdmi_out0_core_initiator_cdc_graycounter0_ce;
assign soc_hdmi_out0_core_initiator_cdc_rdport_adr = soc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary[0];
assign soc_hdmi_out0_core_initiator_cdc_asyncfifo_dout = soc_hdmi_out0_core_initiator_cdc_rdport_dat_r;
always @(*) begin
	soc_hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary <= 2'd0;
	if (soc_hdmi_out0_core_initiator_cdc_graycounter0_ce) begin
		soc_hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary <= (soc_hdmi_out0_core_initiator_cdc_graycounter0_q_binary + 1'd1);
	end else begin
		soc_hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary <= soc_hdmi_out0_core_initiator_cdc_graycounter0_q_binary;
	end
end
assign soc_hdmi_out0_core_initiator_cdc_graycounter0_q_next = (soc_hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary ^ soc_hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary[1]);
always @(*) begin
	soc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary <= 2'd0;
	if (soc_hdmi_out0_core_initiator_cdc_graycounter1_ce) begin
		soc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary <= (soc_hdmi_out0_core_initiator_cdc_graycounter1_q_binary + 1'd1);
	end else begin
		soc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary <= soc_hdmi_out0_core_initiator_cdc_graycounter1_q_binary;
	end
end
assign soc_hdmi_out0_core_initiator_cdc_graycounter1_q_next = (soc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary ^ soc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary[1]);
always @(*) begin
	soc_hdmi_out0_core_timinggenerator_source_valid <= 1'd0;
	soc_hdmi_out0_core_timinggenerator_active <= 1'd0;
	soc_hdmi_out0_core_timinggenerator_source_payload_de <= 1'd0;
	if (soc_hdmi_out0_core_timinggenerator_sink_valid) begin
		soc_hdmi_out0_core_timinggenerator_active <= (soc_hdmi_out0_core_timinggenerator_hactive & soc_hdmi_out0_core_timinggenerator_vactive);
		soc_hdmi_out0_core_timinggenerator_source_valid <= 1'd1;
		if (soc_hdmi_out0_core_timinggenerator_active) begin
			soc_hdmi_out0_core_timinggenerator_source_payload_de <= 1'd1;
		end
	end
end
assign soc_hdmi_out0_core_timinggenerator_sink_ready = (soc_hdmi_out0_core_timinggenerator_source_ready & soc_hdmi_out0_core_timinggenerator_source_last);
assign soc_hdmi_out0_core_dmareader_base = soc_hdmi_out0_core_dmareader_sink_payload_base[31:1];
assign soc_hdmi_out0_core_dmareader_length = soc_hdmi_out0_core_dmareader_sink_payload_length[31:1];
assign soc_hdmi_out0_core_dmareader_sink_sink_payload_address = (soc_hdmi_out0_core_dmareader_base + soc_hdmi_out0_core_dmareader_offset);
assign soc_hdmi_out0_core_dmareader_source_valid = soc_hdmi_out0_core_dmareader_source_source_valid;
assign soc_hdmi_out0_core_dmareader_source_source_ready = soc_hdmi_out0_core_dmareader_source_ready;
assign soc_hdmi_out0_core_dmareader_source_first = soc_hdmi_out0_core_dmareader_source_source_first;
assign soc_hdmi_out0_core_dmareader_source_last = soc_hdmi_out0_core_dmareader_source_source_last;
assign soc_hdmi_out0_core_dmareader_source_payload_data = soc_hdmi_out0_core_dmareader_source_source_payload_data;
assign soc_hdmi_out0_dram_port_litedramport1_cmd_payload_we = 1'd0;
assign soc_hdmi_out0_dram_port_litedramport1_cmd_valid = (soc_hdmi_out0_core_dmareader_sink_sink_valid & soc_hdmi_out0_core_dmareader_request_enable);
assign soc_hdmi_out0_dram_port_litedramport1_cmd_payload_adr = soc_hdmi_out0_core_dmareader_sink_sink_payload_address;
assign soc_hdmi_out0_core_dmareader_sink_sink_ready = (soc_hdmi_out0_dram_port_litedramport1_cmd_ready & soc_hdmi_out0_core_dmareader_request_enable);
assign soc_hdmi_out0_core_dmareader_request_issued = (soc_hdmi_out0_dram_port_litedramport1_cmd_valid & soc_hdmi_out0_dram_port_litedramport1_cmd_ready);
assign soc_hdmi_out0_core_dmareader_request_enable = (soc_hdmi_out0_core_dmareader_rsv_level != 13'd4096);
assign soc_hdmi_out0_core_dmareader_fifo_sink_valid = soc_hdmi_out0_dram_port_litedramport1_rdata_valid;
assign soc_hdmi_out0_dram_port_litedramport1_rdata_ready = soc_hdmi_out0_core_dmareader_fifo_sink_ready;
assign soc_hdmi_out0_core_dmareader_fifo_sink_first = soc_hdmi_out0_dram_port_litedramport1_rdata_first;
assign soc_hdmi_out0_core_dmareader_fifo_sink_last = soc_hdmi_out0_dram_port_litedramport1_rdata_last;
assign soc_hdmi_out0_core_dmareader_fifo_sink_payload_data = soc_hdmi_out0_dram_port_litedramport1_rdata_payload_data;
assign soc_hdmi_out0_core_dmareader_source_source_valid = soc_hdmi_out0_core_dmareader_fifo_source_valid;
assign soc_hdmi_out0_core_dmareader_fifo_source_ready = soc_hdmi_out0_core_dmareader_source_source_ready;
assign soc_hdmi_out0_core_dmareader_source_source_first = soc_hdmi_out0_core_dmareader_fifo_source_first;
assign soc_hdmi_out0_core_dmareader_source_source_last = soc_hdmi_out0_core_dmareader_fifo_source_last;
assign soc_hdmi_out0_core_dmareader_source_source_payload_data = soc_hdmi_out0_core_dmareader_fifo_source_payload_data;
assign soc_hdmi_out0_core_dmareader_data_dequeued = (soc_hdmi_out0_core_dmareader_source_source_valid & soc_hdmi_out0_core_dmareader_source_source_ready);
assign soc_hdmi_out0_core_dmareader_fifo_syncfifo_din = {soc_hdmi_out0_core_dmareader_fifo_fifo_in_last, soc_hdmi_out0_core_dmareader_fifo_fifo_in_first, soc_hdmi_out0_core_dmareader_fifo_fifo_in_payload_data};
assign {soc_hdmi_out0_core_dmareader_fifo_fifo_out_last, soc_hdmi_out0_core_dmareader_fifo_fifo_out_first, soc_hdmi_out0_core_dmareader_fifo_fifo_out_payload_data} = soc_hdmi_out0_core_dmareader_fifo_syncfifo_dout;
assign soc_hdmi_out0_core_dmareader_fifo_sink_ready = soc_hdmi_out0_core_dmareader_fifo_syncfifo_writable;
assign soc_hdmi_out0_core_dmareader_fifo_syncfifo_we = soc_hdmi_out0_core_dmareader_fifo_sink_valid;
assign soc_hdmi_out0_core_dmareader_fifo_fifo_in_first = soc_hdmi_out0_core_dmareader_fifo_sink_first;
assign soc_hdmi_out0_core_dmareader_fifo_fifo_in_last = soc_hdmi_out0_core_dmareader_fifo_sink_last;
assign soc_hdmi_out0_core_dmareader_fifo_fifo_in_payload_data = soc_hdmi_out0_core_dmareader_fifo_sink_payload_data;
assign soc_hdmi_out0_core_dmareader_fifo_source_valid = soc_hdmi_out0_core_dmareader_fifo_readable;
assign soc_hdmi_out0_core_dmareader_fifo_source_first = soc_hdmi_out0_core_dmareader_fifo_fifo_out_first;
assign soc_hdmi_out0_core_dmareader_fifo_source_last = soc_hdmi_out0_core_dmareader_fifo_fifo_out_last;
assign soc_hdmi_out0_core_dmareader_fifo_source_payload_data = soc_hdmi_out0_core_dmareader_fifo_fifo_out_payload_data;
assign soc_hdmi_out0_core_dmareader_fifo_re = soc_hdmi_out0_core_dmareader_fifo_source_ready;
assign soc_hdmi_out0_core_dmareader_fifo_syncfifo_re = (soc_hdmi_out0_core_dmareader_fifo_syncfifo_readable & ((~soc_hdmi_out0_core_dmareader_fifo_readable) | soc_hdmi_out0_core_dmareader_fifo_re));
assign soc_hdmi_out0_core_dmareader_fifo_level1 = (soc_hdmi_out0_core_dmareader_fifo_level0 + soc_hdmi_out0_core_dmareader_fifo_readable);
always @(*) begin
	soc_hdmi_out0_core_dmareader_fifo_wrport_adr <= 12'd0;
	if (soc_hdmi_out0_core_dmareader_fifo_replace) begin
		soc_hdmi_out0_core_dmareader_fifo_wrport_adr <= (soc_hdmi_out0_core_dmareader_fifo_produce - 1'd1);
	end else begin
		soc_hdmi_out0_core_dmareader_fifo_wrport_adr <= soc_hdmi_out0_core_dmareader_fifo_produce;
	end
end
assign soc_hdmi_out0_core_dmareader_fifo_wrport_dat_w = soc_hdmi_out0_core_dmareader_fifo_syncfifo_din;
assign soc_hdmi_out0_core_dmareader_fifo_wrport_we = (soc_hdmi_out0_core_dmareader_fifo_syncfifo_we & (soc_hdmi_out0_core_dmareader_fifo_syncfifo_writable | soc_hdmi_out0_core_dmareader_fifo_replace));
assign soc_hdmi_out0_core_dmareader_fifo_do_read = (soc_hdmi_out0_core_dmareader_fifo_syncfifo_readable & soc_hdmi_out0_core_dmareader_fifo_syncfifo_re);
assign soc_hdmi_out0_core_dmareader_fifo_rdport_adr = soc_hdmi_out0_core_dmareader_fifo_consume;
assign soc_hdmi_out0_core_dmareader_fifo_syncfifo_dout = soc_hdmi_out0_core_dmareader_fifo_rdport_dat_r;
assign soc_hdmi_out0_core_dmareader_fifo_rdport_re = soc_hdmi_out0_core_dmareader_fifo_do_read;
assign soc_hdmi_out0_core_dmareader_fifo_syncfifo_writable = (soc_hdmi_out0_core_dmareader_fifo_level0 != 13'd4096);
assign soc_hdmi_out0_core_dmareader_fifo_syncfifo_readable = (soc_hdmi_out0_core_dmareader_fifo_level0 != 1'd0);
always @(*) begin
	soc_hdmi_out0_core_dmareader_offset_next_value_ce <= 1'd0;
	vns_videoout_next_state <= 1'd0;
	soc_hdmi_out0_core_dmareader_sink_ready <= 1'd0;
	soc_hdmi_out0_dram_port_litedramport1_flush <= 1'd0;
	soc_hdmi_out0_core_dmareader_offset_next_value <= 28'd0;
	soc_hdmi_out0_core_dmareader_sink_sink_valid <= 1'd0;
	vns_videoout_next_state <= vns_videoout_state;
	case (vns_videoout_state)
		1'd1: begin
			soc_hdmi_out0_core_dmareader_sink_sink_valid <= 1'd1;
			if (soc_hdmi_out0_core_dmareader_sink_sink_ready) begin
				soc_hdmi_out0_core_dmareader_offset_next_value <= (soc_hdmi_out0_core_dmareader_offset + 1'd1);
				soc_hdmi_out0_core_dmareader_offset_next_value_ce <= 1'd1;
				if ((soc_hdmi_out0_core_dmareader_offset == (soc_hdmi_out0_core_dmareader_length - 1'd1))) begin
					soc_hdmi_out0_core_dmareader_sink_ready <= 1'd1;
					vns_videoout_next_state <= 1'd0;
				end
			end
		end
		default: begin
			soc_hdmi_out0_core_dmareader_offset_next_value <= 1'd0;
			soc_hdmi_out0_core_dmareader_offset_next_value_ce <= 1'd1;
			if (soc_hdmi_out0_core_dmareader_sink_valid) begin
				vns_videoout_next_state <= 1'd1;
			end else begin
				soc_hdmi_out0_dram_port_litedramport1_flush <= 1'd1;
			end
		end
	endcase
end
assign soc_hdmi_out0_core_o = (soc_hdmi_out0_core_toggle_o ^ soc_hdmi_out0_core_toggle_o_r);
assign soc_hdmi_out0_driver_hdmi_phy_sink_valid = soc_hdmi_out0_driver_sink_sink_valid;
assign soc_hdmi_out0_driver_sink_sink_ready = soc_hdmi_out0_driver_hdmi_phy_sink_ready;
assign soc_hdmi_out0_driver_hdmi_phy_sink_first = soc_hdmi_out0_driver_sink_sink_first;
assign soc_hdmi_out0_driver_hdmi_phy_sink_last = soc_hdmi_out0_driver_sink_sink_last;
assign soc_hdmi_out0_driver_hdmi_phy_sink_payload_r = soc_hdmi_out0_driver_sink_sink_payload_r;
assign soc_hdmi_out0_driver_hdmi_phy_sink_payload_g = soc_hdmi_out0_driver_sink_sink_payload_g;
assign soc_hdmi_out0_driver_hdmi_phy_sink_payload_b = soc_hdmi_out0_driver_sink_sink_payload_b;
assign soc_hdmi_out0_driver_hdmi_phy_sink_param_hsync = soc_hdmi_out0_driver_sink_sink_param_hsync;
assign soc_hdmi_out0_driver_hdmi_phy_sink_param_vsync = soc_hdmi_out0_driver_sink_sink_param_vsync;
assign soc_hdmi_out0_driver_hdmi_phy_sink_param_de = soc_hdmi_out0_driver_sink_sink_param_de;
assign hdmi_out0_pix_rst = (~soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_locked);
assign soc_hdmi_out0_driver_s7hdmioutclocking_data0 = soc_hdmi_out0_driver_s7hdmioutclocking;
assign soc_hdmi_out0_driver_s7hdmioutclocking_data1 = soc_hdmi_out0_driver_s7hdmioutclocking_data0;
assign soc_hdmi_out0_driver_hdmi_phy_sink_ready = 1'd1;
assign soc_hdmi_out0_driver_hdmi_phy_es0_d0 = soc_hdmi_out0_driver_hdmi_phy_sink_payload_b;
assign soc_hdmi_out0_driver_hdmi_phy_es1_d0 = soc_hdmi_out0_driver_hdmi_phy_sink_payload_g;
assign soc_hdmi_out0_driver_hdmi_phy_es2_d0 = soc_hdmi_out0_driver_hdmi_phy_sink_payload_r;
assign soc_hdmi_out0_driver_hdmi_phy_es0_c = {soc_hdmi_out0_driver_hdmi_phy_sink_param_vsync, soc_hdmi_out0_driver_hdmi_phy_sink_param_hsync};
assign soc_hdmi_out0_driver_hdmi_phy_es1_c = 1'd0;
assign soc_hdmi_out0_driver_hdmi_phy_es2_c = 1'd0;
assign soc_hdmi_out0_driver_hdmi_phy_es0_de = soc_hdmi_out0_driver_hdmi_phy_sink_param_de;
assign soc_hdmi_out0_driver_hdmi_phy_es1_de = soc_hdmi_out0_driver_hdmi_phy_sink_param_de;
assign soc_hdmi_out0_driver_hdmi_phy_es2_de = soc_hdmi_out0_driver_hdmi_phy_sink_param_de;
assign soc_hdmi_out0_driver_hdmi_phy_es0_data = soc_hdmi_out0_driver_hdmi_phy_es0_out;
assign soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n = ((soc_hdmi_out0_driver_hdmi_phy_es0_n1d > 3'd4) | ((soc_hdmi_out0_driver_hdmi_phy_es0_n1d == 3'd4) & (~soc_hdmi_out0_driver_hdmi_phy_es0_d1[0])));
assign soc_hdmi_out0_driver_hdmi_phy_es1_data = soc_hdmi_out0_driver_hdmi_phy_es1_out;
assign soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n = ((soc_hdmi_out0_driver_hdmi_phy_es1_n1d > 3'd4) | ((soc_hdmi_out0_driver_hdmi_phy_es1_n1d == 3'd4) & (~soc_hdmi_out0_driver_hdmi_phy_es1_d1[0])));
assign soc_hdmi_out0_driver_hdmi_phy_es2_data = soc_hdmi_out0_driver_hdmi_phy_es2_out;
assign soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n = ((soc_hdmi_out0_driver_hdmi_phy_es2_n1d > 3'd4) | ((soc_hdmi_out0_driver_hdmi_phy_es2_n1d == 3'd4) & (~soc_hdmi_out0_driver_hdmi_phy_es2_d1[0])));
always @(*) begin
	soc_hdmi_out0_resetinserter_cb_fifo_sink_valid <= 1'd0;
	soc_hdmi_out0_resetinserter_cr_fifo_sink_valid <= 1'd0;
	soc_hdmi_out0_resetinserter_sink_sink_ready <= 1'd0;
	soc_hdmi_out0_resetinserter_cb_fifo_sink_payload_data <= 8'd0;
	soc_hdmi_out0_resetinserter_cr_fifo_sink_payload_data <= 8'd0;
	soc_hdmi_out0_resetinserter_y_fifo_sink_payload_data <= 8'd0;
	soc_hdmi_out0_resetinserter_y_fifo_sink_valid <= 1'd0;
	if ((~soc_hdmi_out0_resetinserter_parity_in)) begin
		soc_hdmi_out0_resetinserter_y_fifo_sink_valid <= (soc_hdmi_out0_resetinserter_sink_sink_valid & soc_hdmi_out0_resetinserter_sink_sink_ready);
		soc_hdmi_out0_resetinserter_y_fifo_sink_payload_data <= soc_hdmi_out0_resetinserter_sink_sink_payload_y;
		soc_hdmi_out0_resetinserter_cb_fifo_sink_valid <= (soc_hdmi_out0_resetinserter_sink_sink_valid & soc_hdmi_out0_resetinserter_sink_sink_ready);
		soc_hdmi_out0_resetinserter_cb_fifo_sink_payload_data <= soc_hdmi_out0_resetinserter_sink_sink_payload_cb_cr;
		soc_hdmi_out0_resetinserter_sink_sink_ready <= (soc_hdmi_out0_resetinserter_y_fifo_sink_ready & soc_hdmi_out0_resetinserter_cb_fifo_sink_ready);
	end else begin
		soc_hdmi_out0_resetinserter_y_fifo_sink_valid <= (soc_hdmi_out0_resetinserter_sink_sink_valid & soc_hdmi_out0_resetinserter_sink_sink_ready);
		soc_hdmi_out0_resetinserter_y_fifo_sink_payload_data <= soc_hdmi_out0_resetinserter_sink_sink_payload_y;
		soc_hdmi_out0_resetinserter_cr_fifo_sink_valid <= (soc_hdmi_out0_resetinserter_sink_sink_valid & soc_hdmi_out0_resetinserter_sink_sink_ready);
		soc_hdmi_out0_resetinserter_cr_fifo_sink_payload_data <= soc_hdmi_out0_resetinserter_sink_sink_payload_cb_cr;
		soc_hdmi_out0_resetinserter_sink_sink_ready <= (soc_hdmi_out0_resetinserter_y_fifo_sink_ready & soc_hdmi_out0_resetinserter_cr_fifo_sink_ready);
	end
end
assign soc_hdmi_out0_resetinserter_source_source_valid = ((soc_hdmi_out0_resetinserter_y_fifo_source_valid & soc_hdmi_out0_resetinserter_cb_fifo_source_valid) & soc_hdmi_out0_resetinserter_cr_fifo_source_valid);
assign soc_hdmi_out0_resetinserter_source_source_payload_y = soc_hdmi_out0_resetinserter_y_fifo_source_payload_data;
assign soc_hdmi_out0_resetinserter_source_source_payload_cb = soc_hdmi_out0_resetinserter_cb_fifo_source_payload_data;
assign soc_hdmi_out0_resetinserter_source_source_payload_cr = soc_hdmi_out0_resetinserter_cr_fifo_source_payload_data;
assign soc_hdmi_out0_resetinserter_y_fifo_source_ready = (soc_hdmi_out0_resetinserter_source_source_valid & soc_hdmi_out0_resetinserter_source_source_ready);
assign soc_hdmi_out0_resetinserter_cb_fifo_source_ready = ((soc_hdmi_out0_resetinserter_source_source_valid & soc_hdmi_out0_resetinserter_source_source_ready) & soc_hdmi_out0_resetinserter_parity_out);
assign soc_hdmi_out0_resetinserter_cr_fifo_source_ready = ((soc_hdmi_out0_resetinserter_source_source_valid & soc_hdmi_out0_resetinserter_source_source_ready) & soc_hdmi_out0_resetinserter_parity_out);
assign soc_hdmi_out0_resetinserter_y_fifo_syncfifo_din = {soc_hdmi_out0_resetinserter_y_fifo_fifo_in_last, soc_hdmi_out0_resetinserter_y_fifo_fifo_in_first, soc_hdmi_out0_resetinserter_y_fifo_fifo_in_payload_data};
assign {soc_hdmi_out0_resetinserter_y_fifo_fifo_out_last, soc_hdmi_out0_resetinserter_y_fifo_fifo_out_first, soc_hdmi_out0_resetinserter_y_fifo_fifo_out_payload_data} = soc_hdmi_out0_resetinserter_y_fifo_syncfifo_dout;
assign soc_hdmi_out0_resetinserter_y_fifo_sink_ready = soc_hdmi_out0_resetinserter_y_fifo_syncfifo_writable;
assign soc_hdmi_out0_resetinserter_y_fifo_syncfifo_we = soc_hdmi_out0_resetinserter_y_fifo_sink_valid;
assign soc_hdmi_out0_resetinserter_y_fifo_fifo_in_first = soc_hdmi_out0_resetinserter_y_fifo_sink_first;
assign soc_hdmi_out0_resetinserter_y_fifo_fifo_in_last = soc_hdmi_out0_resetinserter_y_fifo_sink_last;
assign soc_hdmi_out0_resetinserter_y_fifo_fifo_in_payload_data = soc_hdmi_out0_resetinserter_y_fifo_sink_payload_data;
assign soc_hdmi_out0_resetinserter_y_fifo_source_valid = soc_hdmi_out0_resetinserter_y_fifo_syncfifo_readable;
assign soc_hdmi_out0_resetinserter_y_fifo_source_first = soc_hdmi_out0_resetinserter_y_fifo_fifo_out_first;
assign soc_hdmi_out0_resetinserter_y_fifo_source_last = soc_hdmi_out0_resetinserter_y_fifo_fifo_out_last;
assign soc_hdmi_out0_resetinserter_y_fifo_source_payload_data = soc_hdmi_out0_resetinserter_y_fifo_fifo_out_payload_data;
assign soc_hdmi_out0_resetinserter_y_fifo_syncfifo_re = soc_hdmi_out0_resetinserter_y_fifo_source_ready;
always @(*) begin
	soc_hdmi_out0_resetinserter_y_fifo_wrport_adr <= 2'd0;
	if (soc_hdmi_out0_resetinserter_y_fifo_replace) begin
		soc_hdmi_out0_resetinserter_y_fifo_wrport_adr <= (soc_hdmi_out0_resetinserter_y_fifo_produce - 1'd1);
	end else begin
		soc_hdmi_out0_resetinserter_y_fifo_wrport_adr <= soc_hdmi_out0_resetinserter_y_fifo_produce;
	end
end
assign soc_hdmi_out0_resetinserter_y_fifo_wrport_dat_w = soc_hdmi_out0_resetinserter_y_fifo_syncfifo_din;
assign soc_hdmi_out0_resetinserter_y_fifo_wrport_we = (soc_hdmi_out0_resetinserter_y_fifo_syncfifo_we & (soc_hdmi_out0_resetinserter_y_fifo_syncfifo_writable | soc_hdmi_out0_resetinserter_y_fifo_replace));
assign soc_hdmi_out0_resetinserter_y_fifo_do_read = (soc_hdmi_out0_resetinserter_y_fifo_syncfifo_readable & soc_hdmi_out0_resetinserter_y_fifo_syncfifo_re);
assign soc_hdmi_out0_resetinserter_y_fifo_rdport_adr = soc_hdmi_out0_resetinserter_y_fifo_consume;
assign soc_hdmi_out0_resetinserter_y_fifo_syncfifo_dout = soc_hdmi_out0_resetinserter_y_fifo_rdport_dat_r;
assign soc_hdmi_out0_resetinserter_y_fifo_syncfifo_writable = (soc_hdmi_out0_resetinserter_y_fifo_level != 3'd4);
assign soc_hdmi_out0_resetinserter_y_fifo_syncfifo_readable = (soc_hdmi_out0_resetinserter_y_fifo_level != 1'd0);
assign soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_din = {soc_hdmi_out0_resetinserter_cb_fifo_fifo_in_last, soc_hdmi_out0_resetinserter_cb_fifo_fifo_in_first, soc_hdmi_out0_resetinserter_cb_fifo_fifo_in_payload_data};
assign {soc_hdmi_out0_resetinserter_cb_fifo_fifo_out_last, soc_hdmi_out0_resetinserter_cb_fifo_fifo_out_first, soc_hdmi_out0_resetinserter_cb_fifo_fifo_out_payload_data} = soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_dout;
assign soc_hdmi_out0_resetinserter_cb_fifo_sink_ready = soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_writable;
assign soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_we = soc_hdmi_out0_resetinserter_cb_fifo_sink_valid;
assign soc_hdmi_out0_resetinserter_cb_fifo_fifo_in_first = soc_hdmi_out0_resetinserter_cb_fifo_sink_first;
assign soc_hdmi_out0_resetinserter_cb_fifo_fifo_in_last = soc_hdmi_out0_resetinserter_cb_fifo_sink_last;
assign soc_hdmi_out0_resetinserter_cb_fifo_fifo_in_payload_data = soc_hdmi_out0_resetinserter_cb_fifo_sink_payload_data;
assign soc_hdmi_out0_resetinserter_cb_fifo_source_valid = soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_readable;
assign soc_hdmi_out0_resetinserter_cb_fifo_source_first = soc_hdmi_out0_resetinserter_cb_fifo_fifo_out_first;
assign soc_hdmi_out0_resetinserter_cb_fifo_source_last = soc_hdmi_out0_resetinserter_cb_fifo_fifo_out_last;
assign soc_hdmi_out0_resetinserter_cb_fifo_source_payload_data = soc_hdmi_out0_resetinserter_cb_fifo_fifo_out_payload_data;
assign soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_re = soc_hdmi_out0_resetinserter_cb_fifo_source_ready;
always @(*) begin
	soc_hdmi_out0_resetinserter_cb_fifo_wrport_adr <= 2'd0;
	if (soc_hdmi_out0_resetinserter_cb_fifo_replace) begin
		soc_hdmi_out0_resetinserter_cb_fifo_wrport_adr <= (soc_hdmi_out0_resetinserter_cb_fifo_produce - 1'd1);
	end else begin
		soc_hdmi_out0_resetinserter_cb_fifo_wrport_adr <= soc_hdmi_out0_resetinserter_cb_fifo_produce;
	end
end
assign soc_hdmi_out0_resetinserter_cb_fifo_wrport_dat_w = soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_din;
assign soc_hdmi_out0_resetinserter_cb_fifo_wrport_we = (soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_we & (soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_writable | soc_hdmi_out0_resetinserter_cb_fifo_replace));
assign soc_hdmi_out0_resetinserter_cb_fifo_do_read = (soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_readable & soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_re);
assign soc_hdmi_out0_resetinserter_cb_fifo_rdport_adr = soc_hdmi_out0_resetinserter_cb_fifo_consume;
assign soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_dout = soc_hdmi_out0_resetinserter_cb_fifo_rdport_dat_r;
assign soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_writable = (soc_hdmi_out0_resetinserter_cb_fifo_level != 3'd4);
assign soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_readable = (soc_hdmi_out0_resetinserter_cb_fifo_level != 1'd0);
assign soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_din = {soc_hdmi_out0_resetinserter_cr_fifo_fifo_in_last, soc_hdmi_out0_resetinserter_cr_fifo_fifo_in_first, soc_hdmi_out0_resetinserter_cr_fifo_fifo_in_payload_data};
assign {soc_hdmi_out0_resetinserter_cr_fifo_fifo_out_last, soc_hdmi_out0_resetinserter_cr_fifo_fifo_out_first, soc_hdmi_out0_resetinserter_cr_fifo_fifo_out_payload_data} = soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_dout;
assign soc_hdmi_out0_resetinserter_cr_fifo_sink_ready = soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_writable;
assign soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_we = soc_hdmi_out0_resetinserter_cr_fifo_sink_valid;
assign soc_hdmi_out0_resetinserter_cr_fifo_fifo_in_first = soc_hdmi_out0_resetinserter_cr_fifo_sink_first;
assign soc_hdmi_out0_resetinserter_cr_fifo_fifo_in_last = soc_hdmi_out0_resetinserter_cr_fifo_sink_last;
assign soc_hdmi_out0_resetinserter_cr_fifo_fifo_in_payload_data = soc_hdmi_out0_resetinserter_cr_fifo_sink_payload_data;
assign soc_hdmi_out0_resetinserter_cr_fifo_source_valid = soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_readable;
assign soc_hdmi_out0_resetinserter_cr_fifo_source_first = soc_hdmi_out0_resetinserter_cr_fifo_fifo_out_first;
assign soc_hdmi_out0_resetinserter_cr_fifo_source_last = soc_hdmi_out0_resetinserter_cr_fifo_fifo_out_last;
assign soc_hdmi_out0_resetinserter_cr_fifo_source_payload_data = soc_hdmi_out0_resetinserter_cr_fifo_fifo_out_payload_data;
assign soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_re = soc_hdmi_out0_resetinserter_cr_fifo_source_ready;
always @(*) begin
	soc_hdmi_out0_resetinserter_cr_fifo_wrport_adr <= 2'd0;
	if (soc_hdmi_out0_resetinserter_cr_fifo_replace) begin
		soc_hdmi_out0_resetinserter_cr_fifo_wrport_adr <= (soc_hdmi_out0_resetinserter_cr_fifo_produce - 1'd1);
	end else begin
		soc_hdmi_out0_resetinserter_cr_fifo_wrport_adr <= soc_hdmi_out0_resetinserter_cr_fifo_produce;
	end
end
assign soc_hdmi_out0_resetinserter_cr_fifo_wrport_dat_w = soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_din;
assign soc_hdmi_out0_resetinserter_cr_fifo_wrport_we = (soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_we & (soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_writable | soc_hdmi_out0_resetinserter_cr_fifo_replace));
assign soc_hdmi_out0_resetinserter_cr_fifo_do_read = (soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_readable & soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_re);
assign soc_hdmi_out0_resetinserter_cr_fifo_rdport_adr = soc_hdmi_out0_resetinserter_cr_fifo_consume;
assign soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_dout = soc_hdmi_out0_resetinserter_cr_fifo_rdport_dat_r;
assign soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_writable = (soc_hdmi_out0_resetinserter_cr_fifo_level != 3'd4);
assign soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_readable = (soc_hdmi_out0_resetinserter_cr_fifo_level != 1'd0);
assign soc_hdmi_out0_pipe_ce = (soc_hdmi_out0_source_ready | (~soc_hdmi_out0_valid_n3));
assign soc_hdmi_out0_sink_ready = soc_hdmi_out0_pipe_ce;
assign soc_hdmi_out0_source_valid = soc_hdmi_out0_valid_n3;
assign soc_hdmi_out0_busy = ((((1'd0 | soc_hdmi_out0_valid_n0) | soc_hdmi_out0_valid_n1) | soc_hdmi_out0_valid_n2) | soc_hdmi_out0_valid_n3);
assign soc_hdmi_out0_source_first = soc_hdmi_out0_first_n3;
assign soc_hdmi_out0_source_last = soc_hdmi_out0_last_n3;
assign soc_hdmi_out0_ce = soc_hdmi_out0_pipe_ce;
assign soc_hdmi_out0_sink_y = soc_hdmi_out0_sink_payload_y;
assign soc_hdmi_out0_sink_cb = soc_hdmi_out0_sink_payload_cb;
assign soc_hdmi_out0_sink_cr = soc_hdmi_out0_sink_payload_cr;
assign soc_hdmi_out0_source_payload_r = soc_hdmi_out0_source_r;
assign soc_hdmi_out0_source_payload_g = soc_hdmi_out0_source_g;
assign soc_hdmi_out0_source_payload_b = soc_hdmi_out0_source_b;
assign soc_hdmi_out0_source_payload_hsync = soc_hdmi_out0_next_s5;
assign soc_hdmi_out0_source_payload_vsync = soc_hdmi_out0_next_s11;
assign soc_hdmi_out0_source_payload_de = soc_hdmi_out0_next_s17;
assign soc_videosoc_interface0_wb_sdram_adr = vns_comb_rhs_array_muxed38;
assign soc_videosoc_interface0_wb_sdram_dat_w = vns_comb_rhs_array_muxed39;
assign soc_videosoc_interface0_wb_sdram_sel = vns_comb_rhs_array_muxed40;
assign soc_videosoc_interface0_wb_sdram_cyc = vns_comb_rhs_array_muxed41;
assign soc_videosoc_interface0_wb_sdram_stb = vns_comb_rhs_array_muxed42;
assign soc_videosoc_interface0_wb_sdram_we = vns_comb_rhs_array_muxed43;
assign soc_videosoc_interface0_wb_sdram_cti = vns_comb_rhs_array_muxed44;
assign soc_videosoc_interface0_wb_sdram_bte = vns_comb_rhs_array_muxed45;
assign soc_videosoc_interface1_wb_sdram_dat_r = soc_videosoc_interface0_wb_sdram_dat_r;
assign soc_videosoc_interface1_wb_sdram_ack = (soc_videosoc_interface0_wb_sdram_ack & (vns_wb_sdram_con_grant == 1'd0));
assign soc_videosoc_interface1_wb_sdram_err = (soc_videosoc_interface0_wb_sdram_err & (vns_wb_sdram_con_grant == 1'd0));
assign vns_wb_sdram_con_request = {soc_videosoc_interface1_wb_sdram_cyc};
assign vns_wb_sdram_con_grant = 1'd0;
assign vns_videosoc_shared_adr = vns_comb_rhs_array_muxed46;
assign vns_videosoc_shared_dat_w = vns_comb_rhs_array_muxed47;
assign vns_videosoc_shared_sel = vns_comb_rhs_array_muxed48;
assign vns_videosoc_shared_cyc = vns_comb_rhs_array_muxed49;
assign vns_videosoc_shared_stb = vns_comb_rhs_array_muxed50;
assign vns_videosoc_shared_we = vns_comb_rhs_array_muxed51;
assign vns_videosoc_shared_cti = vns_comb_rhs_array_muxed52;
assign vns_videosoc_shared_bte = vns_comb_rhs_array_muxed53;
assign soc_videosoc_videosoc_ibus_dat_r = vns_videosoc_shared_dat_r;
assign soc_videosoc_videosoc_dbus_dat_r = vns_videosoc_shared_dat_r;
assign soc_videosoc_bridge_wishbone_dat_r = vns_videosoc_shared_dat_r;
assign soc_videosoc_videosoc_ibus_ack = (vns_videosoc_shared_ack & (vns_videosoc_grant == 1'd0));
assign soc_videosoc_videosoc_dbus_ack = (vns_videosoc_shared_ack & (vns_videosoc_grant == 1'd1));
assign soc_videosoc_bridge_wishbone_ack = (vns_videosoc_shared_ack & (vns_videosoc_grant == 2'd2));
assign soc_videosoc_videosoc_ibus_err = (vns_videosoc_shared_err & (vns_videosoc_grant == 1'd0));
assign soc_videosoc_videosoc_dbus_err = (vns_videosoc_shared_err & (vns_videosoc_grant == 1'd1));
assign soc_videosoc_bridge_wishbone_err = (vns_videosoc_shared_err & (vns_videosoc_grant == 2'd2));
assign vns_videosoc_request = {soc_videosoc_bridge_wishbone_cyc, soc_videosoc_videosoc_dbus_cyc, soc_videosoc_videosoc_ibus_cyc};
always @(*) begin
	vns_videosoc_slave_sel <= 6'd0;
	vns_videosoc_slave_sel[0] <= (vns_videosoc_shared_adr[28:26] == 1'd0);
	vns_videosoc_slave_sel[1] <= (vns_videosoc_shared_adr[28:26] == 1'd1);
	vns_videosoc_slave_sel[2] <= (vns_videosoc_shared_adr[28:26] == 3'd6);
	vns_videosoc_slave_sel[3] <= (vns_videosoc_shared_adr[28:26] == 3'd4);
	vns_videosoc_slave_sel[4] <= (vns_videosoc_shared_adr[28:26] == 2'd2);
	vns_videosoc_slave_sel[5] <= (vns_videosoc_shared_adr[28:26] == 2'd3);
end
assign soc_videosoc_videosoc_rom_bus_adr = vns_videosoc_shared_adr;
assign soc_videosoc_videosoc_rom_bus_dat_w = vns_videosoc_shared_dat_w;
assign soc_videosoc_videosoc_rom_bus_sel = vns_videosoc_shared_sel;
assign soc_videosoc_videosoc_rom_bus_stb = vns_videosoc_shared_stb;
assign soc_videosoc_videosoc_rom_bus_we = vns_videosoc_shared_we;
assign soc_videosoc_videosoc_rom_bus_cti = vns_videosoc_shared_cti;
assign soc_videosoc_videosoc_rom_bus_bte = vns_videosoc_shared_bte;
assign soc_videosoc_videosoc_sram_bus_adr = vns_videosoc_shared_adr;
assign soc_videosoc_videosoc_sram_bus_dat_w = vns_videosoc_shared_dat_w;
assign soc_videosoc_videosoc_sram_bus_sel = vns_videosoc_shared_sel;
assign soc_videosoc_videosoc_sram_bus_stb = vns_videosoc_shared_stb;
assign soc_videosoc_videosoc_sram_bus_we = vns_videosoc_shared_we;
assign soc_videosoc_videosoc_sram_bus_cti = vns_videosoc_shared_cti;
assign soc_videosoc_videosoc_sram_bus_bte = vns_videosoc_shared_bte;
assign soc_videosoc_videosoc_bus_wishbone_adr = vns_videosoc_shared_adr;
assign soc_videosoc_videosoc_bus_wishbone_dat_w = vns_videosoc_shared_dat_w;
assign soc_videosoc_videosoc_bus_wishbone_sel = vns_videosoc_shared_sel;
assign soc_videosoc_videosoc_bus_wishbone_stb = vns_videosoc_shared_stb;
assign soc_videosoc_videosoc_bus_wishbone_we = vns_videosoc_shared_we;
assign soc_videosoc_videosoc_bus_wishbone_cti = vns_videosoc_shared_cti;
assign soc_videosoc_videosoc_bus_wishbone_bte = vns_videosoc_shared_bte;
assign soc_videosoc_interface1_wb_sdram_adr = vns_videosoc_shared_adr;
assign soc_videosoc_interface1_wb_sdram_dat_w = vns_videosoc_shared_dat_w;
assign soc_videosoc_interface1_wb_sdram_sel = vns_videosoc_shared_sel;
assign soc_videosoc_interface1_wb_sdram_stb = vns_videosoc_shared_stb;
assign soc_videosoc_interface1_wb_sdram_we = vns_videosoc_shared_we;
assign soc_videosoc_interface1_wb_sdram_cti = vns_videosoc_shared_cti;
assign soc_videosoc_interface1_wb_sdram_bte = vns_videosoc_shared_bte;
assign soc_videosoc_bus_adr = vns_videosoc_shared_adr;
assign soc_videosoc_bus_dat_w = vns_videosoc_shared_dat_w;
assign soc_videosoc_bus_sel = vns_videosoc_shared_sel;
assign soc_videosoc_bus_stb = vns_videosoc_shared_stb;
assign soc_videosoc_bus_we = vns_videosoc_shared_we;
assign soc_videosoc_bus_cti = vns_videosoc_shared_cti;
assign soc_videosoc_bus_bte = vns_videosoc_shared_bte;
assign soc_ethmac_bus_adr = vns_videosoc_shared_adr;
assign soc_ethmac_bus_dat_w = vns_videosoc_shared_dat_w;
assign soc_ethmac_bus_sel = vns_videosoc_shared_sel;
assign soc_ethmac_bus_stb = vns_videosoc_shared_stb;
assign soc_ethmac_bus_we = vns_videosoc_shared_we;
assign soc_ethmac_bus_cti = vns_videosoc_shared_cti;
assign soc_ethmac_bus_bte = vns_videosoc_shared_bte;
assign soc_videosoc_videosoc_rom_bus_cyc = (vns_videosoc_shared_cyc & vns_videosoc_slave_sel[0]);
assign soc_videosoc_videosoc_sram_bus_cyc = (vns_videosoc_shared_cyc & vns_videosoc_slave_sel[1]);
assign soc_videosoc_videosoc_bus_wishbone_cyc = (vns_videosoc_shared_cyc & vns_videosoc_slave_sel[2]);
assign soc_videosoc_interface1_wb_sdram_cyc = (vns_videosoc_shared_cyc & vns_videosoc_slave_sel[3]);
assign soc_videosoc_bus_cyc = (vns_videosoc_shared_cyc & vns_videosoc_slave_sel[4]);
assign soc_ethmac_bus_cyc = (vns_videosoc_shared_cyc & vns_videosoc_slave_sel[5]);
assign vns_videosoc_shared_ack = (((((soc_videosoc_videosoc_rom_bus_ack | soc_videosoc_videosoc_sram_bus_ack) | soc_videosoc_videosoc_bus_wishbone_ack) | soc_videosoc_interface1_wb_sdram_ack) | soc_videosoc_bus_ack) | soc_ethmac_bus_ack);
assign vns_videosoc_shared_err = (((((soc_videosoc_videosoc_rom_bus_err | soc_videosoc_videosoc_sram_bus_err) | soc_videosoc_videosoc_bus_wishbone_err) | soc_videosoc_interface1_wb_sdram_err) | soc_videosoc_bus_err) | soc_ethmac_bus_err);
assign vns_videosoc_shared_dat_r = (((((({32{vns_videosoc_slave_sel_r[0]}} & soc_videosoc_videosoc_rom_bus_dat_r) | ({32{vns_videosoc_slave_sel_r[1]}} & soc_videosoc_videosoc_sram_bus_dat_r)) | ({32{vns_videosoc_slave_sel_r[2]}} & soc_videosoc_videosoc_bus_wishbone_dat_r)) | ({32{vns_videosoc_slave_sel_r[3]}} & soc_videosoc_interface1_wb_sdram_dat_r)) | ({32{vns_videosoc_slave_sel_r[4]}} & soc_videosoc_bus_dat_r)) | ({32{vns_videosoc_slave_sel_r[5]}} & soc_ethmac_bus_dat_r));
assign vns_videosoc_csrbank0_sel = (vns_videosoc_interface0_bank_bus_adr[13:9] == 4'd11);
assign vns_videosoc_csrbank0_dly_sel0_r = vns_videosoc_interface0_bank_bus_dat_w[1:0];
assign vns_videosoc_csrbank0_dly_sel0_re = ((vns_videosoc_csrbank0_sel & vns_videosoc_interface0_bank_bus_we) & (vns_videosoc_interface0_bank_bus_adr[1:0] == 1'd0));
assign soc_videosoc_ddrphy_rdly_dq_rst_r = vns_videosoc_interface0_bank_bus_dat_w[0];
assign soc_videosoc_ddrphy_rdly_dq_rst_re = ((vns_videosoc_csrbank0_sel & vns_videosoc_interface0_bank_bus_we) & (vns_videosoc_interface0_bank_bus_adr[1:0] == 1'd1));
assign soc_videosoc_ddrphy_rdly_dq_inc_r = vns_videosoc_interface0_bank_bus_dat_w[0];
assign soc_videosoc_ddrphy_rdly_dq_inc_re = ((vns_videosoc_csrbank0_sel & vns_videosoc_interface0_bank_bus_we) & (vns_videosoc_interface0_bank_bus_adr[1:0] == 2'd2));
assign soc_videosoc_ddrphy_rdly_dq_bitslip_r = vns_videosoc_interface0_bank_bus_dat_w[0];
assign soc_videosoc_ddrphy_rdly_dq_bitslip_re = ((vns_videosoc_csrbank0_sel & vns_videosoc_interface0_bank_bus_we) & (vns_videosoc_interface0_bank_bus_adr[1:0] == 2'd3));
assign soc_videosoc_ddrphy_storage = soc_videosoc_ddrphy_storage_full[1:0];
assign vns_videosoc_csrbank0_dly_sel0_w = soc_videosoc_ddrphy_storage_full[1:0];
assign vns_videosoc_csrbank1_sel = (vns_videosoc_interface1_bank_bus_adr[13:9] == 4'd15);
assign vns_videosoc_csrbank1_sram_writer_slot_r = vns_videosoc_interface1_bank_bus_dat_w[0];
assign vns_videosoc_csrbank1_sram_writer_slot_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 1'd0));
assign vns_videosoc_csrbank1_sram_writer_length3_r = vns_videosoc_interface1_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank1_sram_writer_length3_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 1'd1));
assign vns_videosoc_csrbank1_sram_writer_length2_r = vns_videosoc_interface1_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank1_sram_writer_length2_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 2'd2));
assign vns_videosoc_csrbank1_sram_writer_length1_r = vns_videosoc_interface1_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank1_sram_writer_length1_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 2'd3));
assign vns_videosoc_csrbank1_sram_writer_length0_r = vns_videosoc_interface1_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank1_sram_writer_length0_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 3'd4));
assign soc_ethmac_writer_status_r = vns_videosoc_interface1_bank_bus_dat_w[0];
assign soc_ethmac_writer_status_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 3'd5));
assign soc_ethmac_writer_pending_r = vns_videosoc_interface1_bank_bus_dat_w[0];
assign soc_ethmac_writer_pending_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 3'd6));
assign vns_videosoc_csrbank1_sram_writer_ev_enable0_r = vns_videosoc_interface1_bank_bus_dat_w[0];
assign vns_videosoc_csrbank1_sram_writer_ev_enable0_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 3'd7));
assign soc_ethmac_reader_start_r = vns_videosoc_interface1_bank_bus_dat_w[0];
assign soc_ethmac_reader_start_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 4'd8));
assign vns_videosoc_csrbank1_sram_reader_ready_r = vns_videosoc_interface1_bank_bus_dat_w[0];
assign vns_videosoc_csrbank1_sram_reader_ready_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 4'd9));
assign vns_videosoc_csrbank1_sram_reader_slot0_r = vns_videosoc_interface1_bank_bus_dat_w[0];
assign vns_videosoc_csrbank1_sram_reader_slot0_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 4'd10));
assign vns_videosoc_csrbank1_sram_reader_length1_r = vns_videosoc_interface1_bank_bus_dat_w[2:0];
assign vns_videosoc_csrbank1_sram_reader_length1_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 4'd11));
assign vns_videosoc_csrbank1_sram_reader_length0_r = vns_videosoc_interface1_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank1_sram_reader_length0_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 4'd12));
assign soc_ethmac_reader_eventmanager_status_r = vns_videosoc_interface1_bank_bus_dat_w[0];
assign soc_ethmac_reader_eventmanager_status_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 4'd13));
assign soc_ethmac_reader_eventmanager_pending_r = vns_videosoc_interface1_bank_bus_dat_w[0];
assign soc_ethmac_reader_eventmanager_pending_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 4'd14));
assign vns_videosoc_csrbank1_sram_reader_ev_enable0_r = vns_videosoc_interface1_bank_bus_dat_w[0];
assign vns_videosoc_csrbank1_sram_reader_ev_enable0_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 4'd15));
assign vns_videosoc_csrbank1_preamble_crc_r = vns_videosoc_interface1_bank_bus_dat_w[0];
assign vns_videosoc_csrbank1_preamble_crc_re = ((vns_videosoc_csrbank1_sel & vns_videosoc_interface1_bank_bus_we) & (vns_videosoc_interface1_bank_bus_adr[4:0] == 5'd16));
assign vns_videosoc_csrbank1_sram_writer_slot_w = soc_ethmac_writer_slot_status;
assign vns_videosoc_csrbank1_sram_writer_length3_w = soc_ethmac_writer_length_status[31:24];
assign vns_videosoc_csrbank1_sram_writer_length2_w = soc_ethmac_writer_length_status[23:16];
assign vns_videosoc_csrbank1_sram_writer_length1_w = soc_ethmac_writer_length_status[15:8];
assign vns_videosoc_csrbank1_sram_writer_length0_w = soc_ethmac_writer_length_status[7:0];
assign soc_ethmac_writer_storage = soc_ethmac_writer_storage_full;
assign vns_videosoc_csrbank1_sram_writer_ev_enable0_w = soc_ethmac_writer_storage_full;
assign vns_videosoc_csrbank1_sram_reader_ready_w = soc_ethmac_reader_ready_status;
assign soc_ethmac_reader_slot_storage = soc_ethmac_reader_slot_storage_full;
assign vns_videosoc_csrbank1_sram_reader_slot0_w = soc_ethmac_reader_slot_storage_full;
assign soc_ethmac_reader_length_storage = soc_ethmac_reader_length_storage_full[10:0];
assign vns_videosoc_csrbank1_sram_reader_length1_w = soc_ethmac_reader_length_storage_full[10:8];
assign vns_videosoc_csrbank1_sram_reader_length0_w = soc_ethmac_reader_length_storage_full[7:0];
assign soc_ethmac_reader_eventmanager_storage = soc_ethmac_reader_eventmanager_storage_full;
assign vns_videosoc_csrbank1_sram_reader_ev_enable0_w = soc_ethmac_reader_eventmanager_storage_full;
assign vns_videosoc_csrbank1_preamble_crc_w = soc_ethmac_status;
assign vns_videosoc_csrbank2_sel = (vns_videosoc_interface2_bank_bus_adr[13:9] == 4'd14);
assign vns_videosoc_csrbank2_crg_reset0_r = vns_videosoc_interface2_bank_bus_dat_w[0];
assign vns_videosoc_csrbank2_crg_reset0_re = ((vns_videosoc_csrbank2_sel & vns_videosoc_interface2_bank_bus_we) & (vns_videosoc_interface2_bank_bus_adr[1:0] == 1'd0));
assign vns_videosoc_csrbank2_mdio_w0_r = vns_videosoc_interface2_bank_bus_dat_w[2:0];
assign vns_videosoc_csrbank2_mdio_w0_re = ((vns_videosoc_csrbank2_sel & vns_videosoc_interface2_bank_bus_we) & (vns_videosoc_interface2_bank_bus_adr[1:0] == 1'd1));
assign vns_videosoc_csrbank2_mdio_r_r = vns_videosoc_interface2_bank_bus_dat_w[0];
assign vns_videosoc_csrbank2_mdio_r_re = ((vns_videosoc_csrbank2_sel & vns_videosoc_interface2_bank_bus_we) & (vns_videosoc_interface2_bank_bus_adr[1:0] == 2'd2));
assign soc_ethphy_reset_storage = soc_ethphy_reset_storage_full;
assign vns_videosoc_csrbank2_crg_reset0_w = soc_ethphy_reset_storage_full;
assign soc_ethphy_storage = soc_ethphy_storage_full[2:0];
assign vns_videosoc_csrbank2_mdio_w0_w = soc_ethphy_storage_full[2:0];
assign vns_videosoc_csrbank2_mdio_r_w = soc_ethphy_status;
assign vns_videosoc_sel = (vns_videosoc_sram_bus_adr[13:9] == 5'd19);
always @(*) begin
	vns_videosoc_sram_bus_dat_r <= 8'd0;
	if (vns_videosoc_sel_r) begin
		vns_videosoc_sram_bus_dat_r <= vns_videosoc_dat_r;
	end
end
assign vns_videosoc_we = (vns_videosoc_sel & vns_videosoc_sram_bus_we);
assign vns_videosoc_dat_w = vns_videosoc_sram_bus_dat_w;
assign vns_videosoc_adr = vns_videosoc_sram_bus_adr[6:0];
assign vns_videosoc_csrbank3_sel = (vns_videosoc_interface3_bank_bus_adr[13:9] == 5'd17);
assign vns_videosoc_csrbank3_edid_hpd_notif_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign vns_videosoc_csrbank3_edid_hpd_notif_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 1'd0));
assign vns_videosoc_csrbank3_edid_hpd_en0_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign vns_videosoc_csrbank3_edid_hpd_en0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 1'd1));
assign vns_videosoc_csrbank3_clocking_mmcm_reset0_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign vns_videosoc_csrbank3_clocking_mmcm_reset0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 2'd2));
assign vns_videosoc_csrbank3_clocking_locked_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign vns_videosoc_csrbank3_clocking_locked_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 2'd3));
assign soc_mmcm_read_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign soc_mmcm_read_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 3'd4));
assign soc_mmcm_write_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign soc_mmcm_write_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 3'd5));
assign vns_videosoc_csrbank3_clocking_mmcm_drdy_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign vns_videosoc_csrbank3_clocking_mmcm_drdy_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 3'd6));
assign vns_videosoc_csrbank3_clocking_mmcm_adr0_r = vns_videosoc_interface3_bank_bus_dat_w[6:0];
assign vns_videosoc_csrbank3_clocking_mmcm_adr0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 3'd7));
assign vns_videosoc_csrbank3_clocking_mmcm_dat_w1_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_clocking_mmcm_dat_w1_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 4'd8));
assign vns_videosoc_csrbank3_clocking_mmcm_dat_w0_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_clocking_mmcm_dat_w0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 4'd9));
assign vns_videosoc_csrbank3_clocking_mmcm_dat_r1_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_clocking_mmcm_dat_r1_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 4'd10));
assign vns_videosoc_csrbank3_clocking_mmcm_dat_r0_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_clocking_mmcm_dat_r0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 4'd11));
assign soc_s7datacapture0_dly_ctl_r = vns_videosoc_interface3_bank_bus_dat_w[4:0];
assign soc_s7datacapture0_dly_ctl_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 4'd12));
assign vns_videosoc_csrbank3_data0_cap_phase_r = vns_videosoc_interface3_bank_bus_dat_w[1:0];
assign vns_videosoc_csrbank3_data0_cap_phase_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 4'd13));
assign soc_s7datacapture0_phase_reset_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign soc_s7datacapture0_phase_reset_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 4'd14));
assign vns_videosoc_csrbank3_data0_charsync_char_synced_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign vns_videosoc_csrbank3_data0_charsync_char_synced_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 4'd15));
assign vns_videosoc_csrbank3_data0_charsync_ctl_pos_r = vns_videosoc_interface3_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank3_data0_charsync_ctl_pos_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd16));
assign soc_wer0_update_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign soc_wer0_update_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd17));
assign vns_videosoc_csrbank3_data0_wer_value2_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_data0_wer_value2_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd18));
assign vns_videosoc_csrbank3_data0_wer_value1_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_data0_wer_value1_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd19));
assign vns_videosoc_csrbank3_data0_wer_value0_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_data0_wer_value0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd20));
assign soc_s7datacapture1_dly_ctl_r = vns_videosoc_interface3_bank_bus_dat_w[4:0];
assign soc_s7datacapture1_dly_ctl_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd21));
assign vns_videosoc_csrbank3_data1_cap_phase_r = vns_videosoc_interface3_bank_bus_dat_w[1:0];
assign vns_videosoc_csrbank3_data1_cap_phase_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd22));
assign soc_s7datacapture1_phase_reset_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign soc_s7datacapture1_phase_reset_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd23));
assign vns_videosoc_csrbank3_data1_charsync_char_synced_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign vns_videosoc_csrbank3_data1_charsync_char_synced_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd24));
assign vns_videosoc_csrbank3_data1_charsync_ctl_pos_r = vns_videosoc_interface3_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank3_data1_charsync_ctl_pos_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd25));
assign soc_wer1_update_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign soc_wer1_update_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd26));
assign vns_videosoc_csrbank3_data1_wer_value2_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_data1_wer_value2_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd27));
assign vns_videosoc_csrbank3_data1_wer_value1_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_data1_wer_value1_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd28));
assign vns_videosoc_csrbank3_data1_wer_value0_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_data1_wer_value0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd29));
assign soc_s7datacapture2_dly_ctl_r = vns_videosoc_interface3_bank_bus_dat_w[4:0];
assign soc_s7datacapture2_dly_ctl_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd30));
assign vns_videosoc_csrbank3_data2_cap_phase_r = vns_videosoc_interface3_bank_bus_dat_w[1:0];
assign vns_videosoc_csrbank3_data2_cap_phase_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 5'd31));
assign soc_s7datacapture2_phase_reset_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign soc_s7datacapture2_phase_reset_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd32));
assign vns_videosoc_csrbank3_data2_charsync_char_synced_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign vns_videosoc_csrbank3_data2_charsync_char_synced_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd33));
assign vns_videosoc_csrbank3_data2_charsync_ctl_pos_r = vns_videosoc_interface3_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank3_data2_charsync_ctl_pos_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd34));
assign soc_wer2_update_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign soc_wer2_update_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd35));
assign vns_videosoc_csrbank3_data2_wer_value2_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_data2_wer_value2_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd36));
assign vns_videosoc_csrbank3_data2_wer_value1_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_data2_wer_value1_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd37));
assign vns_videosoc_csrbank3_data2_wer_value0_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_data2_wer_value0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd38));
assign vns_videosoc_csrbank3_chansync_channels_synced_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign vns_videosoc_csrbank3_chansync_channels_synced_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd39));
assign vns_videosoc_csrbank3_resdetection_hres1_r = vns_videosoc_interface3_bank_bus_dat_w[2:0];
assign vns_videosoc_csrbank3_resdetection_hres1_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd40));
assign vns_videosoc_csrbank3_resdetection_hres0_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_resdetection_hres0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd41));
assign vns_videosoc_csrbank3_resdetection_vres1_r = vns_videosoc_interface3_bank_bus_dat_w[2:0];
assign vns_videosoc_csrbank3_resdetection_vres1_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd42));
assign vns_videosoc_csrbank3_resdetection_vres0_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_resdetection_vres0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd43));
assign soc_frame_overflow_r = vns_videosoc_interface3_bank_bus_dat_w[0];
assign soc_frame_overflow_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd44));
assign vns_videosoc_csrbank3_dma_frame_size3_r = vns_videosoc_interface3_bank_bus_dat_w[4:0];
assign vns_videosoc_csrbank3_dma_frame_size3_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd45));
assign vns_videosoc_csrbank3_dma_frame_size2_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_dma_frame_size2_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd46));
assign vns_videosoc_csrbank3_dma_frame_size1_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_dma_frame_size1_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd47));
assign vns_videosoc_csrbank3_dma_frame_size0_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_dma_frame_size0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd48));
assign vns_videosoc_csrbank3_dma_slot0_status0_r = vns_videosoc_interface3_bank_bus_dat_w[1:0];
assign vns_videosoc_csrbank3_dma_slot0_status0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd49));
assign vns_videosoc_csrbank3_dma_slot0_address3_r = vns_videosoc_interface3_bank_bus_dat_w[4:0];
assign vns_videosoc_csrbank3_dma_slot0_address3_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd50));
assign vns_videosoc_csrbank3_dma_slot0_address2_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_dma_slot0_address2_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd51));
assign vns_videosoc_csrbank3_dma_slot0_address1_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_dma_slot0_address1_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd52));
assign vns_videosoc_csrbank3_dma_slot0_address0_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_dma_slot0_address0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd53));
assign vns_videosoc_csrbank3_dma_slot1_status0_r = vns_videosoc_interface3_bank_bus_dat_w[1:0];
assign vns_videosoc_csrbank3_dma_slot1_status0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd54));
assign vns_videosoc_csrbank3_dma_slot1_address3_r = vns_videosoc_interface3_bank_bus_dat_w[4:0];
assign vns_videosoc_csrbank3_dma_slot1_address3_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd55));
assign vns_videosoc_csrbank3_dma_slot1_address2_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_dma_slot1_address2_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd56));
assign vns_videosoc_csrbank3_dma_slot1_address1_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_dma_slot1_address1_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd57));
assign vns_videosoc_csrbank3_dma_slot1_address0_r = vns_videosoc_interface3_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank3_dma_slot1_address0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd58));
assign soc_dma_slot_array_status_r = vns_videosoc_interface3_bank_bus_dat_w[1:0];
assign soc_dma_slot_array_status_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd59));
assign soc_dma_slot_array_pending_r = vns_videosoc_interface3_bank_bus_dat_w[1:0];
assign soc_dma_slot_array_pending_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd60));
assign vns_videosoc_csrbank3_dma_ev_enable0_r = vns_videosoc_interface3_bank_bus_dat_w[1:0];
assign vns_videosoc_csrbank3_dma_ev_enable0_re = ((vns_videosoc_csrbank3_sel & vns_videosoc_interface3_bank_bus_we) & (vns_videosoc_interface3_bank_bus_adr[5:0] == 6'd61));
assign vns_videosoc_csrbank3_edid_hpd_notif_w = soc_edid_status;
assign soc_edid_storage = soc_edid_storage_full;
assign vns_videosoc_csrbank3_edid_hpd_en0_w = soc_edid_storage_full;
assign soc_mmcm_reset_storage = soc_mmcm_reset_storage_full;
assign vns_videosoc_csrbank3_clocking_mmcm_reset0_w = soc_mmcm_reset_storage_full;
assign vns_videosoc_csrbank3_clocking_locked_w = soc_locked_status;
assign vns_videosoc_csrbank3_clocking_mmcm_drdy_w = soc_mmcm_drdy_status;
assign soc_mmcm_adr_storage = soc_mmcm_adr_storage_full[6:0];
assign vns_videosoc_csrbank3_clocking_mmcm_adr0_w = soc_mmcm_adr_storage_full[6:0];
assign soc_mmcm_dat_w_storage = soc_mmcm_dat_w_storage_full[15:0];
assign vns_videosoc_csrbank3_clocking_mmcm_dat_w1_w = soc_mmcm_dat_w_storage_full[15:8];
assign vns_videosoc_csrbank3_clocking_mmcm_dat_w0_w = soc_mmcm_dat_w_storage_full[7:0];
assign vns_videosoc_csrbank3_clocking_mmcm_dat_r1_w = soc_mmcm_dat_r_status[15:8];
assign vns_videosoc_csrbank3_clocking_mmcm_dat_r0_w = soc_mmcm_dat_r_status[7:0];
assign vns_videosoc_csrbank3_data0_cap_phase_w = soc_s7datacapture0_status[1:0];
assign vns_videosoc_csrbank3_data0_charsync_char_synced_w = soc_charsync0_char_synced_status;
assign vns_videosoc_csrbank3_data0_charsync_ctl_pos_w = soc_charsync0_ctl_pos_status[3:0];
assign vns_videosoc_csrbank3_data0_wer_value2_w = soc_wer0_status[23:16];
assign vns_videosoc_csrbank3_data0_wer_value1_w = soc_wer0_status[15:8];
assign vns_videosoc_csrbank3_data0_wer_value0_w = soc_wer0_status[7:0];
assign vns_videosoc_csrbank3_data1_cap_phase_w = soc_s7datacapture1_status[1:0];
assign vns_videosoc_csrbank3_data1_charsync_char_synced_w = soc_charsync1_char_synced_status;
assign vns_videosoc_csrbank3_data1_charsync_ctl_pos_w = soc_charsync1_ctl_pos_status[3:0];
assign vns_videosoc_csrbank3_data1_wer_value2_w = soc_wer1_status[23:16];
assign vns_videosoc_csrbank3_data1_wer_value1_w = soc_wer1_status[15:8];
assign vns_videosoc_csrbank3_data1_wer_value0_w = soc_wer1_status[7:0];
assign vns_videosoc_csrbank3_data2_cap_phase_w = soc_s7datacapture2_status[1:0];
assign vns_videosoc_csrbank3_data2_charsync_char_synced_w = soc_charsync2_char_synced_status;
assign vns_videosoc_csrbank3_data2_charsync_ctl_pos_w = soc_charsync2_ctl_pos_status[3:0];
assign vns_videosoc_csrbank3_data2_wer_value2_w = soc_wer2_status[23:16];
assign vns_videosoc_csrbank3_data2_wer_value1_w = soc_wer2_status[15:8];
assign vns_videosoc_csrbank3_data2_wer_value0_w = soc_wer2_status[7:0];
assign vns_videosoc_csrbank3_chansync_channels_synced_w = soc_chansync_status;
assign vns_videosoc_csrbank3_resdetection_hres1_w = soc_resdetection_hres_status[10:8];
assign vns_videosoc_csrbank3_resdetection_hres0_w = soc_resdetection_hres_status[7:0];
assign vns_videosoc_csrbank3_resdetection_vres1_w = soc_resdetection_vres_status[10:8];
assign vns_videosoc_csrbank3_resdetection_vres0_w = soc_resdetection_vres_status[7:0];
assign soc_dma_frame_size_storage = soc_dma_frame_size_storage_full[28:4];
assign vns_videosoc_csrbank3_dma_frame_size3_w = soc_dma_frame_size_storage_full[28:24];
assign vns_videosoc_csrbank3_dma_frame_size2_w = soc_dma_frame_size_storage_full[23:16];
assign vns_videosoc_csrbank3_dma_frame_size1_w = soc_dma_frame_size_storage_full[15:8];
assign vns_videosoc_csrbank3_dma_frame_size0_w = {soc_dma_frame_size_storage_full[7:4], {4{1'd0}}};
assign soc_dma_slot_array_slot0_status_storage = soc_dma_slot_array_slot0_status_storage_full[1:0];
assign vns_videosoc_csrbank3_dma_slot0_status0_w = soc_dma_slot_array_slot0_status_storage_full[1:0];
assign soc_dma_slot_array_slot0_address_storage = soc_dma_slot_array_slot0_address_storage_full[28:4];
assign vns_videosoc_csrbank3_dma_slot0_address3_w = soc_dma_slot_array_slot0_address_storage_full[28:24];
assign vns_videosoc_csrbank3_dma_slot0_address2_w = soc_dma_slot_array_slot0_address_storage_full[23:16];
assign vns_videosoc_csrbank3_dma_slot0_address1_w = soc_dma_slot_array_slot0_address_storage_full[15:8];
assign vns_videosoc_csrbank3_dma_slot0_address0_w = {soc_dma_slot_array_slot0_address_storage_full[7:4], {4{1'd0}}};
assign soc_dma_slot_array_slot1_status_storage = soc_dma_slot_array_slot1_status_storage_full[1:0];
assign vns_videosoc_csrbank3_dma_slot1_status0_w = soc_dma_slot_array_slot1_status_storage_full[1:0];
assign soc_dma_slot_array_slot1_address_storage = soc_dma_slot_array_slot1_address_storage_full[28:4];
assign vns_videosoc_csrbank3_dma_slot1_address3_w = soc_dma_slot_array_slot1_address_storage_full[28:24];
assign vns_videosoc_csrbank3_dma_slot1_address2_w = soc_dma_slot_array_slot1_address_storage_full[23:16];
assign vns_videosoc_csrbank3_dma_slot1_address1_w = soc_dma_slot_array_slot1_address_storage_full[15:8];
assign vns_videosoc_csrbank3_dma_slot1_address0_w = {soc_dma_slot_array_slot1_address_storage_full[7:4], {4{1'd0}}};
assign soc_dma_slot_array_storage = soc_dma_slot_array_storage_full[1:0];
assign vns_videosoc_csrbank3_dma_ev_enable0_w = soc_dma_slot_array_storage_full[1:0];
assign vns_videosoc_csrbank4_sel = (vns_videosoc_interface4_bank_bus_adr[13:9] == 5'd18);
assign vns_videosoc_csrbank4_value3_r = vns_videosoc_interface4_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank4_value3_re = ((vns_videosoc_csrbank4_sel & vns_videosoc_interface4_bank_bus_we) & (vns_videosoc_interface4_bank_bus_adr[1:0] == 1'd0));
assign vns_videosoc_csrbank4_value2_r = vns_videosoc_interface4_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank4_value2_re = ((vns_videosoc_csrbank4_sel & vns_videosoc_interface4_bank_bus_we) & (vns_videosoc_interface4_bank_bus_adr[1:0] == 1'd1));
assign vns_videosoc_csrbank4_value1_r = vns_videosoc_interface4_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank4_value1_re = ((vns_videosoc_csrbank4_sel & vns_videosoc_interface4_bank_bus_we) & (vns_videosoc_interface4_bank_bus_adr[1:0] == 2'd2));
assign vns_videosoc_csrbank4_value0_r = vns_videosoc_interface4_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank4_value0_re = ((vns_videosoc_csrbank4_sel & vns_videosoc_interface4_bank_bus_we) & (vns_videosoc_interface4_bank_bus_adr[1:0] == 2'd3));
assign vns_videosoc_csrbank4_value3_w = soc_hdmi_in0_freq_status[31:24];
assign vns_videosoc_csrbank4_value2_w = soc_hdmi_in0_freq_status[23:16];
assign vns_videosoc_csrbank4_value1_w = soc_hdmi_in0_freq_status[15:8];
assign vns_videosoc_csrbank4_value0_w = soc_hdmi_in0_freq_status[7:0];
assign vns_videosoc_csrbank5_sel = (vns_videosoc_interface5_bank_bus_adr[13:9] == 5'd16);
assign vns_videosoc_csrbank5_core_underflow_enable0_r = vns_videosoc_interface5_bank_bus_dat_w[0];
assign vns_videosoc_csrbank5_core_underflow_enable0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 1'd0));
assign soc_hdmi_out0_core_underflow_update_underflow_update_r = vns_videosoc_interface5_bank_bus_dat_w[0];
assign soc_hdmi_out0_core_underflow_update_underflow_update_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 1'd1));
assign vns_videosoc_csrbank5_core_underflow_counter3_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_underflow_counter3_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 2'd2));
assign vns_videosoc_csrbank5_core_underflow_counter2_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_underflow_counter2_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 2'd3));
assign vns_videosoc_csrbank5_core_underflow_counter1_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_underflow_counter1_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 3'd4));
assign vns_videosoc_csrbank5_core_underflow_counter0_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_underflow_counter0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 3'd5));
assign vns_videosoc_csrbank5_core_initiator_enable0_r = vns_videosoc_interface5_bank_bus_dat_w[0];
assign vns_videosoc_csrbank5_core_initiator_enable0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 3'd6));
assign vns_videosoc_csrbank5_core_initiator_hres1_r = vns_videosoc_interface5_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank5_core_initiator_hres1_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 3'd7));
assign vns_videosoc_csrbank5_core_initiator_hres0_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_hres0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 4'd8));
assign vns_videosoc_csrbank5_core_initiator_hsync_start1_r = vns_videosoc_interface5_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank5_core_initiator_hsync_start1_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 4'd9));
assign vns_videosoc_csrbank5_core_initiator_hsync_start0_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_hsync_start0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 4'd10));
assign vns_videosoc_csrbank5_core_initiator_hsync_end1_r = vns_videosoc_interface5_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank5_core_initiator_hsync_end1_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 4'd11));
assign vns_videosoc_csrbank5_core_initiator_hsync_end0_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_hsync_end0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 4'd12));
assign vns_videosoc_csrbank5_core_initiator_hscan1_r = vns_videosoc_interface5_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank5_core_initiator_hscan1_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 4'd13));
assign vns_videosoc_csrbank5_core_initiator_hscan0_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_hscan0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 4'd14));
assign vns_videosoc_csrbank5_core_initiator_vres1_r = vns_videosoc_interface5_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank5_core_initiator_vres1_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 4'd15));
assign vns_videosoc_csrbank5_core_initiator_vres0_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_vres0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd16));
assign vns_videosoc_csrbank5_core_initiator_vsync_start1_r = vns_videosoc_interface5_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank5_core_initiator_vsync_start1_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd17));
assign vns_videosoc_csrbank5_core_initiator_vsync_start0_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_vsync_start0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd18));
assign vns_videosoc_csrbank5_core_initiator_vsync_end1_r = vns_videosoc_interface5_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank5_core_initiator_vsync_end1_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd19));
assign vns_videosoc_csrbank5_core_initiator_vsync_end0_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_vsync_end0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd20));
assign vns_videosoc_csrbank5_core_initiator_vscan1_r = vns_videosoc_interface5_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank5_core_initiator_vscan1_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd21));
assign vns_videosoc_csrbank5_core_initiator_vscan0_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_vscan0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd22));
assign vns_videosoc_csrbank5_core_initiator_base3_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_base3_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd23));
assign vns_videosoc_csrbank5_core_initiator_base2_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_base2_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd24));
assign vns_videosoc_csrbank5_core_initiator_base1_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_base1_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd25));
assign vns_videosoc_csrbank5_core_initiator_base0_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_base0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd26));
assign vns_videosoc_csrbank5_core_initiator_length3_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_length3_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd27));
assign vns_videosoc_csrbank5_core_initiator_length2_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_length2_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd28));
assign vns_videosoc_csrbank5_core_initiator_length1_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_length1_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd29));
assign vns_videosoc_csrbank5_core_initiator_length0_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_core_initiator_length0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd30));
assign vns_videosoc_csrbank5_driver_clocking_mmcm_reset0_r = vns_videosoc_interface5_bank_bus_dat_w[0];
assign vns_videosoc_csrbank5_driver_clocking_mmcm_reset0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 5'd31));
assign soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_read_r = vns_videosoc_interface5_bank_bus_dat_w[0];
assign soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_read_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 6'd32));
assign soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_write_r = vns_videosoc_interface5_bank_bus_dat_w[0];
assign soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_write_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 6'd33));
assign vns_videosoc_csrbank5_driver_clocking_mmcm_drdy_r = vns_videosoc_interface5_bank_bus_dat_w[0];
assign vns_videosoc_csrbank5_driver_clocking_mmcm_drdy_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 6'd34));
assign vns_videosoc_csrbank5_driver_clocking_mmcm_adr0_r = vns_videosoc_interface5_bank_bus_dat_w[6:0];
assign vns_videosoc_csrbank5_driver_clocking_mmcm_adr0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 6'd35));
assign vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w1_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w1_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 6'd36));
assign vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w0_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 6'd37));
assign vns_videosoc_csrbank5_driver_clocking_mmcm_dat_r1_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_driver_clocking_mmcm_dat_r1_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 6'd38));
assign vns_videosoc_csrbank5_driver_clocking_mmcm_dat_r0_r = vns_videosoc_interface5_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank5_driver_clocking_mmcm_dat_r0_re = ((vns_videosoc_csrbank5_sel & vns_videosoc_interface5_bank_bus_we) & (vns_videosoc_interface5_bank_bus_adr[5:0] == 6'd39));
assign soc_hdmi_out0_core_underflow_enable_storage = soc_hdmi_out0_core_underflow_enable_storage_full;
assign vns_videosoc_csrbank5_core_underflow_enable0_w = soc_hdmi_out0_core_underflow_enable_storage_full;
assign vns_videosoc_csrbank5_core_underflow_counter3_w = soc_hdmi_out0_core_underflow_counter_status[31:24];
assign vns_videosoc_csrbank5_core_underflow_counter2_w = soc_hdmi_out0_core_underflow_counter_status[23:16];
assign vns_videosoc_csrbank5_core_underflow_counter1_w = soc_hdmi_out0_core_underflow_counter_status[15:8];
assign vns_videosoc_csrbank5_core_underflow_counter0_w = soc_hdmi_out0_core_underflow_counter_status[7:0];
assign soc_hdmi_out0_core_initiator_enable_storage = soc_hdmi_out0_core_initiator_enable_storage_full;
assign vns_videosoc_csrbank5_core_initiator_enable0_w = soc_hdmi_out0_core_initiator_enable_storage_full;
assign soc_hdmi_out0_core_initiator_csrstorage0_storage = soc_hdmi_out0_core_initiator_csrstorage0_storage_full[11:0];
assign vns_videosoc_csrbank5_core_initiator_hres1_w = soc_hdmi_out0_core_initiator_csrstorage0_storage_full[11:8];
assign vns_videosoc_csrbank5_core_initiator_hres0_w = soc_hdmi_out0_core_initiator_csrstorage0_storage_full[7:0];
assign soc_hdmi_out0_core_initiator_csrstorage1_storage = soc_hdmi_out0_core_initiator_csrstorage1_storage_full[11:0];
assign vns_videosoc_csrbank5_core_initiator_hsync_start1_w = soc_hdmi_out0_core_initiator_csrstorage1_storage_full[11:8];
assign vns_videosoc_csrbank5_core_initiator_hsync_start0_w = soc_hdmi_out0_core_initiator_csrstorage1_storage_full[7:0];
assign soc_hdmi_out0_core_initiator_csrstorage2_storage = soc_hdmi_out0_core_initiator_csrstorage2_storage_full[11:0];
assign vns_videosoc_csrbank5_core_initiator_hsync_end1_w = soc_hdmi_out0_core_initiator_csrstorage2_storage_full[11:8];
assign vns_videosoc_csrbank5_core_initiator_hsync_end0_w = soc_hdmi_out0_core_initiator_csrstorage2_storage_full[7:0];
assign soc_hdmi_out0_core_initiator_csrstorage3_storage = soc_hdmi_out0_core_initiator_csrstorage3_storage_full[11:0];
assign vns_videosoc_csrbank5_core_initiator_hscan1_w = soc_hdmi_out0_core_initiator_csrstorage3_storage_full[11:8];
assign vns_videosoc_csrbank5_core_initiator_hscan0_w = soc_hdmi_out0_core_initiator_csrstorage3_storage_full[7:0];
assign soc_hdmi_out0_core_initiator_csrstorage4_storage = soc_hdmi_out0_core_initiator_csrstorage4_storage_full[11:0];
assign vns_videosoc_csrbank5_core_initiator_vres1_w = soc_hdmi_out0_core_initiator_csrstorage4_storage_full[11:8];
assign vns_videosoc_csrbank5_core_initiator_vres0_w = soc_hdmi_out0_core_initiator_csrstorage4_storage_full[7:0];
assign soc_hdmi_out0_core_initiator_csrstorage5_storage = soc_hdmi_out0_core_initiator_csrstorage5_storage_full[11:0];
assign vns_videosoc_csrbank5_core_initiator_vsync_start1_w = soc_hdmi_out0_core_initiator_csrstorage5_storage_full[11:8];
assign vns_videosoc_csrbank5_core_initiator_vsync_start0_w = soc_hdmi_out0_core_initiator_csrstorage5_storage_full[7:0];
assign soc_hdmi_out0_core_initiator_csrstorage6_storage = soc_hdmi_out0_core_initiator_csrstorage6_storage_full[11:0];
assign vns_videosoc_csrbank5_core_initiator_vsync_end1_w = soc_hdmi_out0_core_initiator_csrstorage6_storage_full[11:8];
assign vns_videosoc_csrbank5_core_initiator_vsync_end0_w = soc_hdmi_out0_core_initiator_csrstorage6_storage_full[7:0];
assign soc_hdmi_out0_core_initiator_csrstorage7_storage = soc_hdmi_out0_core_initiator_csrstorage7_storage_full[11:0];
assign vns_videosoc_csrbank5_core_initiator_vscan1_w = soc_hdmi_out0_core_initiator_csrstorage7_storage_full[11:8];
assign vns_videosoc_csrbank5_core_initiator_vscan0_w = soc_hdmi_out0_core_initiator_csrstorage7_storage_full[7:0];
assign soc_hdmi_out0_core_initiator_csrstorage8_storage = soc_hdmi_out0_core_initiator_csrstorage8_storage_full[31:0];
assign vns_videosoc_csrbank5_core_initiator_base3_w = soc_hdmi_out0_core_initiator_csrstorage8_storage_full[31:24];
assign vns_videosoc_csrbank5_core_initiator_base2_w = soc_hdmi_out0_core_initiator_csrstorage8_storage_full[23:16];
assign vns_videosoc_csrbank5_core_initiator_base1_w = soc_hdmi_out0_core_initiator_csrstorage8_storage_full[15:8];
assign vns_videosoc_csrbank5_core_initiator_base0_w = soc_hdmi_out0_core_initiator_csrstorage8_storage_full[7:0];
assign soc_hdmi_out0_core_initiator_csrstorage9_storage = soc_hdmi_out0_core_initiator_csrstorage9_storage_full[31:0];
assign vns_videosoc_csrbank5_core_initiator_length3_w = soc_hdmi_out0_core_initiator_csrstorage9_storage_full[31:24];
assign vns_videosoc_csrbank5_core_initiator_length2_w = soc_hdmi_out0_core_initiator_csrstorage9_storage_full[23:16];
assign vns_videosoc_csrbank5_core_initiator_length1_w = soc_hdmi_out0_core_initiator_csrstorage9_storage_full[15:8];
assign vns_videosoc_csrbank5_core_initiator_length0_w = soc_hdmi_out0_core_initiator_csrstorage9_storage_full[7:0];
assign soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage = soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage_full;
assign vns_videosoc_csrbank5_driver_clocking_mmcm_reset0_w = soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage_full;
assign vns_videosoc_csrbank5_driver_clocking_mmcm_drdy_w = soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy_status;
assign soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage = soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage_full[6:0];
assign vns_videosoc_csrbank5_driver_clocking_mmcm_adr0_w = soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage_full[6:0];
assign soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage = soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage_full[15:0];
assign vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w1_w = soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage_full[15:8];
assign vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w0_w = soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage_full[7:0];
assign vns_videosoc_csrbank5_driver_clocking_mmcm_dat_r1_w = soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_r_status[15:8];
assign vns_videosoc_csrbank5_driver_clocking_mmcm_dat_r0_w = soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_r_status[7:0];
assign vns_videosoc_csrbank6_sel = (vns_videosoc_interface6_bank_bus_adr[13:9] == 4'd12);
assign vns_videosoc_csrbank6_dna_id7_r = vns_videosoc_interface6_bank_bus_dat_w[0];
assign vns_videosoc_csrbank6_dna_id7_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 1'd0));
assign vns_videosoc_csrbank6_dna_id6_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_dna_id6_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 1'd1));
assign vns_videosoc_csrbank6_dna_id5_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_dna_id5_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 2'd2));
assign vns_videosoc_csrbank6_dna_id4_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_dna_id4_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 2'd3));
assign vns_videosoc_csrbank6_dna_id3_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_dna_id3_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 3'd4));
assign vns_videosoc_csrbank6_dna_id2_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_dna_id2_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 3'd5));
assign vns_videosoc_csrbank6_dna_id1_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_dna_id1_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 3'd6));
assign vns_videosoc_csrbank6_dna_id0_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_dna_id0_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 3'd7));
assign vns_videosoc_csrbank6_git_commit19_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit19_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 4'd8));
assign vns_videosoc_csrbank6_git_commit18_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit18_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 4'd9));
assign vns_videosoc_csrbank6_git_commit17_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit17_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 4'd10));
assign vns_videosoc_csrbank6_git_commit16_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit16_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 4'd11));
assign vns_videosoc_csrbank6_git_commit15_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit15_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 4'd12));
assign vns_videosoc_csrbank6_git_commit14_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit14_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 4'd13));
assign vns_videosoc_csrbank6_git_commit13_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit13_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 4'd14));
assign vns_videosoc_csrbank6_git_commit12_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit12_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 4'd15));
assign vns_videosoc_csrbank6_git_commit11_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit11_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd16));
assign vns_videosoc_csrbank6_git_commit10_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit10_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd17));
assign vns_videosoc_csrbank6_git_commit9_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit9_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd18));
assign vns_videosoc_csrbank6_git_commit8_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit8_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd19));
assign vns_videosoc_csrbank6_git_commit7_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit7_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd20));
assign vns_videosoc_csrbank6_git_commit6_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit6_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd21));
assign vns_videosoc_csrbank6_git_commit5_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit5_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd22));
assign vns_videosoc_csrbank6_git_commit4_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit4_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd23));
assign vns_videosoc_csrbank6_git_commit3_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit3_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd24));
assign vns_videosoc_csrbank6_git_commit2_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit2_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd25));
assign vns_videosoc_csrbank6_git_commit1_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit1_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd26));
assign vns_videosoc_csrbank6_git_commit0_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_git_commit0_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd27));
assign vns_videosoc_csrbank6_platform_platform7_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_platform7_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd28));
assign vns_videosoc_csrbank6_platform_platform6_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_platform6_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd29));
assign vns_videosoc_csrbank6_platform_platform5_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_platform5_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd30));
assign vns_videosoc_csrbank6_platform_platform4_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_platform4_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 5'd31));
assign vns_videosoc_csrbank6_platform_platform3_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_platform3_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd32));
assign vns_videosoc_csrbank6_platform_platform2_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_platform2_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd33));
assign vns_videosoc_csrbank6_platform_platform1_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_platform1_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd34));
assign vns_videosoc_csrbank6_platform_platform0_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_platform0_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd35));
assign vns_videosoc_csrbank6_platform_target7_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_target7_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd36));
assign vns_videosoc_csrbank6_platform_target6_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_target6_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd37));
assign vns_videosoc_csrbank6_platform_target5_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_target5_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd38));
assign vns_videosoc_csrbank6_platform_target4_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_target4_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd39));
assign vns_videosoc_csrbank6_platform_target3_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_target3_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd40));
assign vns_videosoc_csrbank6_platform_target2_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_target2_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd41));
assign vns_videosoc_csrbank6_platform_target1_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_target1_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd42));
assign vns_videosoc_csrbank6_platform_target0_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_platform_target0_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd43));
assign vns_videosoc_csrbank6_xadc_temperature1_r = vns_videosoc_interface6_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank6_xadc_temperature1_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd44));
assign vns_videosoc_csrbank6_xadc_temperature0_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_xadc_temperature0_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd45));
assign vns_videosoc_csrbank6_xadc_vccint1_r = vns_videosoc_interface6_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank6_xadc_vccint1_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd46));
assign vns_videosoc_csrbank6_xadc_vccint0_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_xadc_vccint0_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd47));
assign vns_videosoc_csrbank6_xadc_vccaux1_r = vns_videosoc_interface6_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank6_xadc_vccaux1_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd48));
assign vns_videosoc_csrbank6_xadc_vccaux0_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_xadc_vccaux0_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd49));
assign vns_videosoc_csrbank6_xadc_vccbram1_r = vns_videosoc_interface6_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank6_xadc_vccbram1_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd50));
assign vns_videosoc_csrbank6_xadc_vccbram0_r = vns_videosoc_interface6_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank6_xadc_vccbram0_re = ((vns_videosoc_csrbank6_sel & vns_videosoc_interface6_bank_bus_we) & (vns_videosoc_interface6_bank_bus_adr[5:0] == 6'd51));
assign vns_videosoc_csrbank6_dna_id7_w = soc_videosoc_info_dna_status[56];
assign vns_videosoc_csrbank6_dna_id6_w = soc_videosoc_info_dna_status[55:48];
assign vns_videosoc_csrbank6_dna_id5_w = soc_videosoc_info_dna_status[47:40];
assign vns_videosoc_csrbank6_dna_id4_w = soc_videosoc_info_dna_status[39:32];
assign vns_videosoc_csrbank6_dna_id3_w = soc_videosoc_info_dna_status[31:24];
assign vns_videosoc_csrbank6_dna_id2_w = soc_videosoc_info_dna_status[23:16];
assign vns_videosoc_csrbank6_dna_id1_w = soc_videosoc_info_dna_status[15:8];
assign vns_videosoc_csrbank6_dna_id0_w = soc_videosoc_info_dna_status[7:0];
assign vns_videosoc_csrbank6_git_commit19_w = soc_videosoc_info_git_status[159:152];
assign vns_videosoc_csrbank6_git_commit18_w = soc_videosoc_info_git_status[151:144];
assign vns_videosoc_csrbank6_git_commit17_w = soc_videosoc_info_git_status[143:136];
assign vns_videosoc_csrbank6_git_commit16_w = soc_videosoc_info_git_status[135:128];
assign vns_videosoc_csrbank6_git_commit15_w = soc_videosoc_info_git_status[127:120];
assign vns_videosoc_csrbank6_git_commit14_w = soc_videosoc_info_git_status[119:112];
assign vns_videosoc_csrbank6_git_commit13_w = soc_videosoc_info_git_status[111:104];
assign vns_videosoc_csrbank6_git_commit12_w = soc_videosoc_info_git_status[103:96];
assign vns_videosoc_csrbank6_git_commit11_w = soc_videosoc_info_git_status[95:88];
assign vns_videosoc_csrbank6_git_commit10_w = soc_videosoc_info_git_status[87:80];
assign vns_videosoc_csrbank6_git_commit9_w = soc_videosoc_info_git_status[79:72];
assign vns_videosoc_csrbank6_git_commit8_w = soc_videosoc_info_git_status[71:64];
assign vns_videosoc_csrbank6_git_commit7_w = soc_videosoc_info_git_status[63:56];
assign vns_videosoc_csrbank6_git_commit6_w = soc_videosoc_info_git_status[55:48];
assign vns_videosoc_csrbank6_git_commit5_w = soc_videosoc_info_git_status[47:40];
assign vns_videosoc_csrbank6_git_commit4_w = soc_videosoc_info_git_status[39:32];
assign vns_videosoc_csrbank6_git_commit3_w = soc_videosoc_info_git_status[31:24];
assign vns_videosoc_csrbank6_git_commit2_w = soc_videosoc_info_git_status[23:16];
assign vns_videosoc_csrbank6_git_commit1_w = soc_videosoc_info_git_status[15:8];
assign vns_videosoc_csrbank6_git_commit0_w = soc_videosoc_info_git_status[7:0];
assign vns_videosoc_csrbank6_platform_platform7_w = soc_videosoc_info_platform_status[63:56];
assign vns_videosoc_csrbank6_platform_platform6_w = soc_videosoc_info_platform_status[55:48];
assign vns_videosoc_csrbank6_platform_platform5_w = soc_videosoc_info_platform_status[47:40];
assign vns_videosoc_csrbank6_platform_platform4_w = soc_videosoc_info_platform_status[39:32];
assign vns_videosoc_csrbank6_platform_platform3_w = soc_videosoc_info_platform_status[31:24];
assign vns_videosoc_csrbank6_platform_platform2_w = soc_videosoc_info_platform_status[23:16];
assign vns_videosoc_csrbank6_platform_platform1_w = soc_videosoc_info_platform_status[15:8];
assign vns_videosoc_csrbank6_platform_platform0_w = soc_videosoc_info_platform_status[7:0];
assign vns_videosoc_csrbank6_platform_target7_w = soc_videosoc_info_target_status[63:56];
assign vns_videosoc_csrbank6_platform_target6_w = soc_videosoc_info_target_status[55:48];
assign vns_videosoc_csrbank6_platform_target5_w = soc_videosoc_info_target_status[47:40];
assign vns_videosoc_csrbank6_platform_target4_w = soc_videosoc_info_target_status[39:32];
assign vns_videosoc_csrbank6_platform_target3_w = soc_videosoc_info_target_status[31:24];
assign vns_videosoc_csrbank6_platform_target2_w = soc_videosoc_info_target_status[23:16];
assign vns_videosoc_csrbank6_platform_target1_w = soc_videosoc_info_target_status[15:8];
assign vns_videosoc_csrbank6_platform_target0_w = soc_videosoc_info_target_status[7:0];
assign vns_videosoc_csrbank6_xadc_temperature1_w = soc_videosoc_info_temperature_status[11:8];
assign vns_videosoc_csrbank6_xadc_temperature0_w = soc_videosoc_info_temperature_status[7:0];
assign vns_videosoc_csrbank6_xadc_vccint1_w = soc_videosoc_info_vccint_status[11:8];
assign vns_videosoc_csrbank6_xadc_vccint0_w = soc_videosoc_info_vccint_status[7:0];
assign vns_videosoc_csrbank6_xadc_vccaux1_w = soc_videosoc_info_vccaux_status[11:8];
assign vns_videosoc_csrbank6_xadc_vccaux0_w = soc_videosoc_info_vccaux_status[7:0];
assign vns_videosoc_csrbank6_xadc_vccbram1_w = soc_videosoc_info_vccbram_status[11:8];
assign vns_videosoc_csrbank6_xadc_vccbram0_w = soc_videosoc_info_vccbram_status[7:0];
assign vns_videosoc_csrbank7_sel = (vns_videosoc_interface7_bank_bus_adr[13:9] == 4'd13);
assign soc_videosoc_oled_spimaster_ctrl_r = vns_videosoc_interface7_bank_bus_dat_w[0];
assign soc_videosoc_oled_spimaster_ctrl_re = ((vns_videosoc_csrbank7_sel & vns_videosoc_interface7_bank_bus_we) & (vns_videosoc_interface7_bank_bus_adr[2:0] == 1'd0));
assign vns_videosoc_csrbank7_spi_length0_r = vns_videosoc_interface7_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank7_spi_length0_re = ((vns_videosoc_csrbank7_sel & vns_videosoc_interface7_bank_bus_we) & (vns_videosoc_interface7_bank_bus_adr[2:0] == 1'd1));
assign vns_videosoc_csrbank7_spi_status_r = vns_videosoc_interface7_bank_bus_dat_w[0];
assign vns_videosoc_csrbank7_spi_status_re = ((vns_videosoc_csrbank7_sel & vns_videosoc_interface7_bank_bus_we) & (vns_videosoc_interface7_bank_bus_adr[2:0] == 2'd2));
assign vns_videosoc_csrbank7_spi_mosi0_r = vns_videosoc_interface7_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank7_spi_mosi0_re = ((vns_videosoc_csrbank7_sel & vns_videosoc_interface7_bank_bus_we) & (vns_videosoc_interface7_bank_bus_adr[2:0] == 2'd3));
assign vns_videosoc_csrbank7_gpio_out0_r = vns_videosoc_interface7_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank7_gpio_out0_re = ((vns_videosoc_csrbank7_sel & vns_videosoc_interface7_bank_bus_we) & (vns_videosoc_interface7_bank_bus_adr[2:0] == 3'd4));
assign soc_videosoc_oled_spimaster_length_storage = soc_videosoc_oled_spimaster_length_storage_full[7:0];
assign vns_videosoc_csrbank7_spi_length0_w = soc_videosoc_oled_spimaster_length_storage_full[7:0];
assign vns_videosoc_csrbank7_spi_status_w = soc_videosoc_oled_spimaster_status;
assign soc_videosoc_oled_spimaster_mosi_storage = soc_videosoc_oled_spimaster_mosi_storage_full[7:0];
assign vns_videosoc_csrbank7_spi_mosi0_w = soc_videosoc_oled_spimaster_mosi_storage_full[7:0];
assign soc_videosoc_oled_storage = soc_videosoc_oled_storage_full[3:0];
assign vns_videosoc_csrbank7_gpio_out0_w = soc_videosoc_oled_storage_full[3:0];
assign vns_videosoc_csrbank8_sel = (vns_videosoc_interface8_bank_bus_adr[13:9] == 4'd8);
assign vns_videosoc_csrbank8_dfii_control0_r = vns_videosoc_interface8_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank8_dfii_control0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 1'd0));
assign vns_videosoc_csrbank8_dfii_pi0_command0_r = vns_videosoc_interface8_bank_bus_dat_w[5:0];
assign vns_videosoc_csrbank8_dfii_pi0_command0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 1'd1));
assign soc_videosoc_sdram_phaseinjector0_command_issue_r = vns_videosoc_interface8_bank_bus_dat_w[0];
assign soc_videosoc_sdram_phaseinjector0_command_issue_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 2'd2));
assign vns_videosoc_csrbank8_dfii_pi0_address1_r = vns_videosoc_interface8_bank_bus_dat_w[6:0];
assign vns_videosoc_csrbank8_dfii_pi0_address1_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 2'd3));
assign vns_videosoc_csrbank8_dfii_pi0_address0_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi0_address0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 3'd4));
assign vns_videosoc_csrbank8_dfii_pi0_baddress0_r = vns_videosoc_interface8_bank_bus_dat_w[2:0];
assign vns_videosoc_csrbank8_dfii_pi0_baddress0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 3'd5));
assign vns_videosoc_csrbank8_dfii_pi0_wrdata3_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi0_wrdata3_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 3'd6));
assign vns_videosoc_csrbank8_dfii_pi0_wrdata2_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi0_wrdata2_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 3'd7));
assign vns_videosoc_csrbank8_dfii_pi0_wrdata1_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi0_wrdata1_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 4'd8));
assign vns_videosoc_csrbank8_dfii_pi0_wrdata0_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi0_wrdata0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 4'd9));
assign vns_videosoc_csrbank8_dfii_pi0_rddata3_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi0_rddata3_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 4'd10));
assign vns_videosoc_csrbank8_dfii_pi0_rddata2_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi0_rddata2_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 4'd11));
assign vns_videosoc_csrbank8_dfii_pi0_rddata1_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi0_rddata1_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 4'd12));
assign vns_videosoc_csrbank8_dfii_pi0_rddata0_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi0_rddata0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 4'd13));
assign vns_videosoc_csrbank8_dfii_pi1_command0_r = vns_videosoc_interface8_bank_bus_dat_w[5:0];
assign vns_videosoc_csrbank8_dfii_pi1_command0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 4'd14));
assign soc_videosoc_sdram_phaseinjector1_command_issue_r = vns_videosoc_interface8_bank_bus_dat_w[0];
assign soc_videosoc_sdram_phaseinjector1_command_issue_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 4'd15));
assign vns_videosoc_csrbank8_dfii_pi1_address1_r = vns_videosoc_interface8_bank_bus_dat_w[6:0];
assign vns_videosoc_csrbank8_dfii_pi1_address1_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd16));
assign vns_videosoc_csrbank8_dfii_pi1_address0_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi1_address0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd17));
assign vns_videosoc_csrbank8_dfii_pi1_baddress0_r = vns_videosoc_interface8_bank_bus_dat_w[2:0];
assign vns_videosoc_csrbank8_dfii_pi1_baddress0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd18));
assign vns_videosoc_csrbank8_dfii_pi1_wrdata3_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi1_wrdata3_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd19));
assign vns_videosoc_csrbank8_dfii_pi1_wrdata2_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi1_wrdata2_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd20));
assign vns_videosoc_csrbank8_dfii_pi1_wrdata1_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi1_wrdata1_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd21));
assign vns_videosoc_csrbank8_dfii_pi1_wrdata0_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi1_wrdata0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd22));
assign vns_videosoc_csrbank8_dfii_pi1_rddata3_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi1_rddata3_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd23));
assign vns_videosoc_csrbank8_dfii_pi1_rddata2_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi1_rddata2_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd24));
assign vns_videosoc_csrbank8_dfii_pi1_rddata1_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi1_rddata1_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd25));
assign vns_videosoc_csrbank8_dfii_pi1_rddata0_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi1_rddata0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd26));
assign vns_videosoc_csrbank8_dfii_pi2_command0_r = vns_videosoc_interface8_bank_bus_dat_w[5:0];
assign vns_videosoc_csrbank8_dfii_pi2_command0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd27));
assign soc_videosoc_sdram_phaseinjector2_command_issue_r = vns_videosoc_interface8_bank_bus_dat_w[0];
assign soc_videosoc_sdram_phaseinjector2_command_issue_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd28));
assign vns_videosoc_csrbank8_dfii_pi2_address1_r = vns_videosoc_interface8_bank_bus_dat_w[6:0];
assign vns_videosoc_csrbank8_dfii_pi2_address1_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd29));
assign vns_videosoc_csrbank8_dfii_pi2_address0_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi2_address0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd30));
assign vns_videosoc_csrbank8_dfii_pi2_baddress0_r = vns_videosoc_interface8_bank_bus_dat_w[2:0];
assign vns_videosoc_csrbank8_dfii_pi2_baddress0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 5'd31));
assign vns_videosoc_csrbank8_dfii_pi2_wrdata3_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi2_wrdata3_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd32));
assign vns_videosoc_csrbank8_dfii_pi2_wrdata2_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi2_wrdata2_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd33));
assign vns_videosoc_csrbank8_dfii_pi2_wrdata1_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi2_wrdata1_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd34));
assign vns_videosoc_csrbank8_dfii_pi2_wrdata0_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi2_wrdata0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd35));
assign vns_videosoc_csrbank8_dfii_pi2_rddata3_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi2_rddata3_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd36));
assign vns_videosoc_csrbank8_dfii_pi2_rddata2_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi2_rddata2_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd37));
assign vns_videosoc_csrbank8_dfii_pi2_rddata1_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi2_rddata1_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd38));
assign vns_videosoc_csrbank8_dfii_pi2_rddata0_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi2_rddata0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd39));
assign vns_videosoc_csrbank8_dfii_pi3_command0_r = vns_videosoc_interface8_bank_bus_dat_w[5:0];
assign vns_videosoc_csrbank8_dfii_pi3_command0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd40));
assign soc_videosoc_sdram_phaseinjector3_command_issue_r = vns_videosoc_interface8_bank_bus_dat_w[0];
assign soc_videosoc_sdram_phaseinjector3_command_issue_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd41));
assign vns_videosoc_csrbank8_dfii_pi3_address1_r = vns_videosoc_interface8_bank_bus_dat_w[6:0];
assign vns_videosoc_csrbank8_dfii_pi3_address1_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd42));
assign vns_videosoc_csrbank8_dfii_pi3_address0_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi3_address0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd43));
assign vns_videosoc_csrbank8_dfii_pi3_baddress0_r = vns_videosoc_interface8_bank_bus_dat_w[2:0];
assign vns_videosoc_csrbank8_dfii_pi3_baddress0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd44));
assign vns_videosoc_csrbank8_dfii_pi3_wrdata3_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi3_wrdata3_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd45));
assign vns_videosoc_csrbank8_dfii_pi3_wrdata2_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi3_wrdata2_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd46));
assign vns_videosoc_csrbank8_dfii_pi3_wrdata1_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi3_wrdata1_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd47));
assign vns_videosoc_csrbank8_dfii_pi3_wrdata0_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi3_wrdata0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd48));
assign vns_videosoc_csrbank8_dfii_pi3_rddata3_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi3_rddata3_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd49));
assign vns_videosoc_csrbank8_dfii_pi3_rddata2_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi3_rddata2_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd50));
assign vns_videosoc_csrbank8_dfii_pi3_rddata1_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi3_rddata1_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd51));
assign vns_videosoc_csrbank8_dfii_pi3_rddata0_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_dfii_pi3_rddata0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd52));
assign soc_videosoc_sdram_bandwidth_update_r = vns_videosoc_interface8_bank_bus_dat_w[0];
assign soc_videosoc_sdram_bandwidth_update_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd53));
assign vns_videosoc_csrbank8_controller_bandwidth_nreads2_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_controller_bandwidth_nreads2_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd54));
assign vns_videosoc_csrbank8_controller_bandwidth_nreads1_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_controller_bandwidth_nreads1_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd55));
assign vns_videosoc_csrbank8_controller_bandwidth_nreads0_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_controller_bandwidth_nreads0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd56));
assign vns_videosoc_csrbank8_controller_bandwidth_nwrites2_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_controller_bandwidth_nwrites2_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd57));
assign vns_videosoc_csrbank8_controller_bandwidth_nwrites1_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_controller_bandwidth_nwrites1_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd58));
assign vns_videosoc_csrbank8_controller_bandwidth_nwrites0_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_controller_bandwidth_nwrites0_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd59));
assign vns_videosoc_csrbank8_controller_bandwidth_data_width_r = vns_videosoc_interface8_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank8_controller_bandwidth_data_width_re = ((vns_videosoc_csrbank8_sel & vns_videosoc_interface8_bank_bus_we) & (vns_videosoc_interface8_bank_bus_adr[5:0] == 6'd60));
assign soc_videosoc_sdram_storage = soc_videosoc_sdram_storage_full[3:0];
assign vns_videosoc_csrbank8_dfii_control0_w = soc_videosoc_sdram_storage_full[3:0];
assign soc_videosoc_sdram_phaseinjector0_command_storage = soc_videosoc_sdram_phaseinjector0_command_storage_full[5:0];
assign vns_videosoc_csrbank8_dfii_pi0_command0_w = soc_videosoc_sdram_phaseinjector0_command_storage_full[5:0];
assign soc_videosoc_sdram_phaseinjector0_address_storage = soc_videosoc_sdram_phaseinjector0_address_storage_full[14:0];
assign vns_videosoc_csrbank8_dfii_pi0_address1_w = soc_videosoc_sdram_phaseinjector0_address_storage_full[14:8];
assign vns_videosoc_csrbank8_dfii_pi0_address0_w = soc_videosoc_sdram_phaseinjector0_address_storage_full[7:0];
assign soc_videosoc_sdram_phaseinjector0_baddress_storage = soc_videosoc_sdram_phaseinjector0_baddress_storage_full[2:0];
assign vns_videosoc_csrbank8_dfii_pi0_baddress0_w = soc_videosoc_sdram_phaseinjector0_baddress_storage_full[2:0];
assign soc_videosoc_sdram_phaseinjector0_wrdata_storage = soc_videosoc_sdram_phaseinjector0_wrdata_storage_full[31:0];
assign vns_videosoc_csrbank8_dfii_pi0_wrdata3_w = soc_videosoc_sdram_phaseinjector0_wrdata_storage_full[31:24];
assign vns_videosoc_csrbank8_dfii_pi0_wrdata2_w = soc_videosoc_sdram_phaseinjector0_wrdata_storage_full[23:16];
assign vns_videosoc_csrbank8_dfii_pi0_wrdata1_w = soc_videosoc_sdram_phaseinjector0_wrdata_storage_full[15:8];
assign vns_videosoc_csrbank8_dfii_pi0_wrdata0_w = soc_videosoc_sdram_phaseinjector0_wrdata_storage_full[7:0];
assign vns_videosoc_csrbank8_dfii_pi0_rddata3_w = soc_videosoc_sdram_phaseinjector0_status[31:24];
assign vns_videosoc_csrbank8_dfii_pi0_rddata2_w = soc_videosoc_sdram_phaseinjector0_status[23:16];
assign vns_videosoc_csrbank8_dfii_pi0_rddata1_w = soc_videosoc_sdram_phaseinjector0_status[15:8];
assign vns_videosoc_csrbank8_dfii_pi0_rddata0_w = soc_videosoc_sdram_phaseinjector0_status[7:0];
assign soc_videosoc_sdram_phaseinjector1_command_storage = soc_videosoc_sdram_phaseinjector1_command_storage_full[5:0];
assign vns_videosoc_csrbank8_dfii_pi1_command0_w = soc_videosoc_sdram_phaseinjector1_command_storage_full[5:0];
assign soc_videosoc_sdram_phaseinjector1_address_storage = soc_videosoc_sdram_phaseinjector1_address_storage_full[14:0];
assign vns_videosoc_csrbank8_dfii_pi1_address1_w = soc_videosoc_sdram_phaseinjector1_address_storage_full[14:8];
assign vns_videosoc_csrbank8_dfii_pi1_address0_w = soc_videosoc_sdram_phaseinjector1_address_storage_full[7:0];
assign soc_videosoc_sdram_phaseinjector1_baddress_storage = soc_videosoc_sdram_phaseinjector1_baddress_storage_full[2:0];
assign vns_videosoc_csrbank8_dfii_pi1_baddress0_w = soc_videosoc_sdram_phaseinjector1_baddress_storage_full[2:0];
assign soc_videosoc_sdram_phaseinjector1_wrdata_storage = soc_videosoc_sdram_phaseinjector1_wrdata_storage_full[31:0];
assign vns_videosoc_csrbank8_dfii_pi1_wrdata3_w = soc_videosoc_sdram_phaseinjector1_wrdata_storage_full[31:24];
assign vns_videosoc_csrbank8_dfii_pi1_wrdata2_w = soc_videosoc_sdram_phaseinjector1_wrdata_storage_full[23:16];
assign vns_videosoc_csrbank8_dfii_pi1_wrdata1_w = soc_videosoc_sdram_phaseinjector1_wrdata_storage_full[15:8];
assign vns_videosoc_csrbank8_dfii_pi1_wrdata0_w = soc_videosoc_sdram_phaseinjector1_wrdata_storage_full[7:0];
assign vns_videosoc_csrbank8_dfii_pi1_rddata3_w = soc_videosoc_sdram_phaseinjector1_status[31:24];
assign vns_videosoc_csrbank8_dfii_pi1_rddata2_w = soc_videosoc_sdram_phaseinjector1_status[23:16];
assign vns_videosoc_csrbank8_dfii_pi1_rddata1_w = soc_videosoc_sdram_phaseinjector1_status[15:8];
assign vns_videosoc_csrbank8_dfii_pi1_rddata0_w = soc_videosoc_sdram_phaseinjector1_status[7:0];
assign soc_videosoc_sdram_phaseinjector2_command_storage = soc_videosoc_sdram_phaseinjector2_command_storage_full[5:0];
assign vns_videosoc_csrbank8_dfii_pi2_command0_w = soc_videosoc_sdram_phaseinjector2_command_storage_full[5:0];
assign soc_videosoc_sdram_phaseinjector2_address_storage = soc_videosoc_sdram_phaseinjector2_address_storage_full[14:0];
assign vns_videosoc_csrbank8_dfii_pi2_address1_w = soc_videosoc_sdram_phaseinjector2_address_storage_full[14:8];
assign vns_videosoc_csrbank8_dfii_pi2_address0_w = soc_videosoc_sdram_phaseinjector2_address_storage_full[7:0];
assign soc_videosoc_sdram_phaseinjector2_baddress_storage = soc_videosoc_sdram_phaseinjector2_baddress_storage_full[2:0];
assign vns_videosoc_csrbank8_dfii_pi2_baddress0_w = soc_videosoc_sdram_phaseinjector2_baddress_storage_full[2:0];
assign soc_videosoc_sdram_phaseinjector2_wrdata_storage = soc_videosoc_sdram_phaseinjector2_wrdata_storage_full[31:0];
assign vns_videosoc_csrbank8_dfii_pi2_wrdata3_w = soc_videosoc_sdram_phaseinjector2_wrdata_storage_full[31:24];
assign vns_videosoc_csrbank8_dfii_pi2_wrdata2_w = soc_videosoc_sdram_phaseinjector2_wrdata_storage_full[23:16];
assign vns_videosoc_csrbank8_dfii_pi2_wrdata1_w = soc_videosoc_sdram_phaseinjector2_wrdata_storage_full[15:8];
assign vns_videosoc_csrbank8_dfii_pi2_wrdata0_w = soc_videosoc_sdram_phaseinjector2_wrdata_storage_full[7:0];
assign vns_videosoc_csrbank8_dfii_pi2_rddata3_w = soc_videosoc_sdram_phaseinjector2_status[31:24];
assign vns_videosoc_csrbank8_dfii_pi2_rddata2_w = soc_videosoc_sdram_phaseinjector2_status[23:16];
assign vns_videosoc_csrbank8_dfii_pi2_rddata1_w = soc_videosoc_sdram_phaseinjector2_status[15:8];
assign vns_videosoc_csrbank8_dfii_pi2_rddata0_w = soc_videosoc_sdram_phaseinjector2_status[7:0];
assign soc_videosoc_sdram_phaseinjector3_command_storage = soc_videosoc_sdram_phaseinjector3_command_storage_full[5:0];
assign vns_videosoc_csrbank8_dfii_pi3_command0_w = soc_videosoc_sdram_phaseinjector3_command_storage_full[5:0];
assign soc_videosoc_sdram_phaseinjector3_address_storage = soc_videosoc_sdram_phaseinjector3_address_storage_full[14:0];
assign vns_videosoc_csrbank8_dfii_pi3_address1_w = soc_videosoc_sdram_phaseinjector3_address_storage_full[14:8];
assign vns_videosoc_csrbank8_dfii_pi3_address0_w = soc_videosoc_sdram_phaseinjector3_address_storage_full[7:0];
assign soc_videosoc_sdram_phaseinjector3_baddress_storage = soc_videosoc_sdram_phaseinjector3_baddress_storage_full[2:0];
assign vns_videosoc_csrbank8_dfii_pi3_baddress0_w = soc_videosoc_sdram_phaseinjector3_baddress_storage_full[2:0];
assign soc_videosoc_sdram_phaseinjector3_wrdata_storage = soc_videosoc_sdram_phaseinjector3_wrdata_storage_full[31:0];
assign vns_videosoc_csrbank8_dfii_pi3_wrdata3_w = soc_videosoc_sdram_phaseinjector3_wrdata_storage_full[31:24];
assign vns_videosoc_csrbank8_dfii_pi3_wrdata2_w = soc_videosoc_sdram_phaseinjector3_wrdata_storage_full[23:16];
assign vns_videosoc_csrbank8_dfii_pi3_wrdata1_w = soc_videosoc_sdram_phaseinjector3_wrdata_storage_full[15:8];
assign vns_videosoc_csrbank8_dfii_pi3_wrdata0_w = soc_videosoc_sdram_phaseinjector3_wrdata_storage_full[7:0];
assign vns_videosoc_csrbank8_dfii_pi3_rddata3_w = soc_videosoc_sdram_phaseinjector3_status[31:24];
assign vns_videosoc_csrbank8_dfii_pi3_rddata2_w = soc_videosoc_sdram_phaseinjector3_status[23:16];
assign vns_videosoc_csrbank8_dfii_pi3_rddata1_w = soc_videosoc_sdram_phaseinjector3_status[15:8];
assign vns_videosoc_csrbank8_dfii_pi3_rddata0_w = soc_videosoc_sdram_phaseinjector3_status[7:0];
assign vns_videosoc_csrbank8_controller_bandwidth_nreads2_w = soc_videosoc_sdram_bandwidth_nreads_status[23:16];
assign vns_videosoc_csrbank8_controller_bandwidth_nreads1_w = soc_videosoc_sdram_bandwidth_nreads_status[15:8];
assign vns_videosoc_csrbank8_controller_bandwidth_nreads0_w = soc_videosoc_sdram_bandwidth_nreads_status[7:0];
assign vns_videosoc_csrbank8_controller_bandwidth_nwrites2_w = soc_videosoc_sdram_bandwidth_nwrites_status[23:16];
assign vns_videosoc_csrbank8_controller_bandwidth_nwrites1_w = soc_videosoc_sdram_bandwidth_nwrites_status[15:8];
assign vns_videosoc_csrbank8_controller_bandwidth_nwrites0_w = soc_videosoc_sdram_bandwidth_nwrites_status[7:0];
assign vns_videosoc_csrbank8_controller_bandwidth_data_width_w = soc_videosoc_sdram_bandwidth_data_width_status[7:0];
assign vns_videosoc_csrbank9_sel = (vns_videosoc_interface9_bank_bus_adr[13:9] == 4'd10);
assign vns_videosoc_csrbank9_bitbang0_r = vns_videosoc_interface9_bank_bus_dat_w[3:0];
assign vns_videosoc_csrbank9_bitbang0_re = ((vns_videosoc_csrbank9_sel & vns_videosoc_interface9_bank_bus_we) & (vns_videosoc_interface9_bank_bus_adr[1:0] == 1'd0));
assign vns_videosoc_csrbank9_miso_r = vns_videosoc_interface9_bank_bus_dat_w[0];
assign vns_videosoc_csrbank9_miso_re = ((vns_videosoc_csrbank9_sel & vns_videosoc_interface9_bank_bus_we) & (vns_videosoc_interface9_bank_bus_adr[1:0] == 1'd1));
assign vns_videosoc_csrbank9_bitbang_en0_r = vns_videosoc_interface9_bank_bus_dat_w[0];
assign vns_videosoc_csrbank9_bitbang_en0_re = ((vns_videosoc_csrbank9_sel & vns_videosoc_interface9_bank_bus_we) & (vns_videosoc_interface9_bank_bus_adr[1:0] == 2'd2));
assign soc_videosoc_bitbang_storage = soc_videosoc_bitbang_storage_full[3:0];
assign vns_videosoc_csrbank9_bitbang0_w = soc_videosoc_bitbang_storage_full[3:0];
assign vns_videosoc_csrbank9_miso_w = soc_videosoc_miso_status;
assign soc_videosoc_bitbang_en_storage = soc_videosoc_bitbang_en_storage_full;
assign vns_videosoc_csrbank9_bitbang_en0_w = soc_videosoc_bitbang_en_storage_full;
assign vns_videosoc_csrbank10_sel = (vns_videosoc_interface10_bank_bus_adr[13:9] == 3'd4);
assign vns_videosoc_csrbank10_load3_r = vns_videosoc_interface10_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank10_load3_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 1'd0));
assign vns_videosoc_csrbank10_load2_r = vns_videosoc_interface10_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank10_load2_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 1'd1));
assign vns_videosoc_csrbank10_load1_r = vns_videosoc_interface10_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank10_load1_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 2'd2));
assign vns_videosoc_csrbank10_load0_r = vns_videosoc_interface10_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank10_load0_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 2'd3));
assign vns_videosoc_csrbank10_reload3_r = vns_videosoc_interface10_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank10_reload3_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 3'd4));
assign vns_videosoc_csrbank10_reload2_r = vns_videosoc_interface10_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank10_reload2_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 3'd5));
assign vns_videosoc_csrbank10_reload1_r = vns_videosoc_interface10_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank10_reload1_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 3'd6));
assign vns_videosoc_csrbank10_reload0_r = vns_videosoc_interface10_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank10_reload0_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 3'd7));
assign vns_videosoc_csrbank10_en0_r = vns_videosoc_interface10_bank_bus_dat_w[0];
assign vns_videosoc_csrbank10_en0_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 4'd8));
assign soc_videosoc_videosoc_update_value_r = vns_videosoc_interface10_bank_bus_dat_w[0];
assign soc_videosoc_videosoc_update_value_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 4'd9));
assign vns_videosoc_csrbank10_value3_r = vns_videosoc_interface10_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank10_value3_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 4'd10));
assign vns_videosoc_csrbank10_value2_r = vns_videosoc_interface10_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank10_value2_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 4'd11));
assign vns_videosoc_csrbank10_value1_r = vns_videosoc_interface10_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank10_value1_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 4'd12));
assign vns_videosoc_csrbank10_value0_r = vns_videosoc_interface10_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank10_value0_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 4'd13));
assign soc_videosoc_videosoc_eventmanager_status_r = vns_videosoc_interface10_bank_bus_dat_w[0];
assign soc_videosoc_videosoc_eventmanager_status_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 4'd14));
assign soc_videosoc_videosoc_eventmanager_pending_r = vns_videosoc_interface10_bank_bus_dat_w[0];
assign soc_videosoc_videosoc_eventmanager_pending_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 4'd15));
assign vns_videosoc_csrbank10_ev_enable0_r = vns_videosoc_interface10_bank_bus_dat_w[0];
assign vns_videosoc_csrbank10_ev_enable0_re = ((vns_videosoc_csrbank10_sel & vns_videosoc_interface10_bank_bus_we) & (vns_videosoc_interface10_bank_bus_adr[4:0] == 5'd16));
assign soc_videosoc_videosoc_load_storage = soc_videosoc_videosoc_load_storage_full[31:0];
assign vns_videosoc_csrbank10_load3_w = soc_videosoc_videosoc_load_storage_full[31:24];
assign vns_videosoc_csrbank10_load2_w = soc_videosoc_videosoc_load_storage_full[23:16];
assign vns_videosoc_csrbank10_load1_w = soc_videosoc_videosoc_load_storage_full[15:8];
assign vns_videosoc_csrbank10_load0_w = soc_videosoc_videosoc_load_storage_full[7:0];
assign soc_videosoc_videosoc_reload_storage = soc_videosoc_videosoc_reload_storage_full[31:0];
assign vns_videosoc_csrbank10_reload3_w = soc_videosoc_videosoc_reload_storage_full[31:24];
assign vns_videosoc_csrbank10_reload2_w = soc_videosoc_videosoc_reload_storage_full[23:16];
assign vns_videosoc_csrbank10_reload1_w = soc_videosoc_videosoc_reload_storage_full[15:8];
assign vns_videosoc_csrbank10_reload0_w = soc_videosoc_videosoc_reload_storage_full[7:0];
assign soc_videosoc_videosoc_en_storage = soc_videosoc_videosoc_en_storage_full;
assign vns_videosoc_csrbank10_en0_w = soc_videosoc_videosoc_en_storage_full;
assign vns_videosoc_csrbank10_value3_w = soc_videosoc_videosoc_value_status[31:24];
assign vns_videosoc_csrbank10_value2_w = soc_videosoc_videosoc_value_status[23:16];
assign vns_videosoc_csrbank10_value1_w = soc_videosoc_videosoc_value_status[15:8];
assign vns_videosoc_csrbank10_value0_w = soc_videosoc_videosoc_value_status[7:0];
assign soc_videosoc_videosoc_eventmanager_storage = soc_videosoc_videosoc_eventmanager_storage_full;
assign vns_videosoc_csrbank10_ev_enable0_w = soc_videosoc_videosoc_eventmanager_storage_full;
assign vns_videosoc_csrbank11_sel = (vns_videosoc_interface11_bank_bus_adr[13:9] == 2'd2);
assign soc_videosoc_uart_rxtx_r = vns_videosoc_interface11_bank_bus_dat_w[7:0];
assign soc_videosoc_uart_rxtx_re = ((vns_videosoc_csrbank11_sel & vns_videosoc_interface11_bank_bus_we) & (vns_videosoc_interface11_bank_bus_adr[2:0] == 1'd0));
assign vns_videosoc_csrbank11_txfull_r = vns_videosoc_interface11_bank_bus_dat_w[0];
assign vns_videosoc_csrbank11_txfull_re = ((vns_videosoc_csrbank11_sel & vns_videosoc_interface11_bank_bus_we) & (vns_videosoc_interface11_bank_bus_adr[2:0] == 1'd1));
assign vns_videosoc_csrbank11_rxempty_r = vns_videosoc_interface11_bank_bus_dat_w[0];
assign vns_videosoc_csrbank11_rxempty_re = ((vns_videosoc_csrbank11_sel & vns_videosoc_interface11_bank_bus_we) & (vns_videosoc_interface11_bank_bus_adr[2:0] == 2'd2));
assign soc_videosoc_uart_status_r = vns_videosoc_interface11_bank_bus_dat_w[1:0];
assign soc_videosoc_uart_status_re = ((vns_videosoc_csrbank11_sel & vns_videosoc_interface11_bank_bus_we) & (vns_videosoc_interface11_bank_bus_adr[2:0] == 2'd3));
assign soc_videosoc_uart_pending_r = vns_videosoc_interface11_bank_bus_dat_w[1:0];
assign soc_videosoc_uart_pending_re = ((vns_videosoc_csrbank11_sel & vns_videosoc_interface11_bank_bus_we) & (vns_videosoc_interface11_bank_bus_adr[2:0] == 3'd4));
assign vns_videosoc_csrbank11_ev_enable0_r = vns_videosoc_interface11_bank_bus_dat_w[1:0];
assign vns_videosoc_csrbank11_ev_enable0_re = ((vns_videosoc_csrbank11_sel & vns_videosoc_interface11_bank_bus_we) & (vns_videosoc_interface11_bank_bus_adr[2:0] == 3'd5));
assign vns_videosoc_csrbank11_txfull_w = soc_videosoc_uart_txfull_status;
assign vns_videosoc_csrbank11_rxempty_w = soc_videosoc_uart_rxempty_status;
assign soc_videosoc_uart_storage = soc_videosoc_uart_storage_full[1:0];
assign vns_videosoc_csrbank11_ev_enable0_w = soc_videosoc_uart_storage_full[1:0];
assign vns_videosoc_csrbank12_sel = (vns_videosoc_interface12_bank_bus_adr[13:9] == 1'd1);
assign vns_videosoc_csrbank12_tuning_word3_r = vns_videosoc_interface12_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank12_tuning_word3_re = ((vns_videosoc_csrbank12_sel & vns_videosoc_interface12_bank_bus_we) & (vns_videosoc_interface12_bank_bus_adr[1:0] == 1'd0));
assign vns_videosoc_csrbank12_tuning_word2_r = vns_videosoc_interface12_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank12_tuning_word2_re = ((vns_videosoc_csrbank12_sel & vns_videosoc_interface12_bank_bus_we) & (vns_videosoc_interface12_bank_bus_adr[1:0] == 1'd1));
assign vns_videosoc_csrbank12_tuning_word1_r = vns_videosoc_interface12_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank12_tuning_word1_re = ((vns_videosoc_csrbank12_sel & vns_videosoc_interface12_bank_bus_we) & (vns_videosoc_interface12_bank_bus_adr[1:0] == 2'd2));
assign vns_videosoc_csrbank12_tuning_word0_r = vns_videosoc_interface12_bank_bus_dat_w[7:0];
assign vns_videosoc_csrbank12_tuning_word0_re = ((vns_videosoc_csrbank12_sel & vns_videosoc_interface12_bank_bus_we) & (vns_videosoc_interface12_bank_bus_adr[1:0] == 2'd3));
assign soc_videosoc_uart_phy_storage = soc_videosoc_uart_phy_storage_full[31:0];
assign vns_videosoc_csrbank12_tuning_word3_w = soc_videosoc_uart_phy_storage_full[31:24];
assign vns_videosoc_csrbank12_tuning_word2_w = soc_videosoc_uart_phy_storage_full[23:16];
assign vns_videosoc_csrbank12_tuning_word1_w = soc_videosoc_uart_phy_storage_full[15:8];
assign vns_videosoc_csrbank12_tuning_word0_w = soc_videosoc_uart_phy_storage_full[7:0];
assign vns_videosoc_interface0_bank_bus_adr = soc_videosoc_videosoc_interface_adr;
assign vns_videosoc_interface1_bank_bus_adr = soc_videosoc_videosoc_interface_adr;
assign vns_videosoc_interface2_bank_bus_adr = soc_videosoc_videosoc_interface_adr;
assign vns_videosoc_interface3_bank_bus_adr = soc_videosoc_videosoc_interface_adr;
assign vns_videosoc_interface4_bank_bus_adr = soc_videosoc_videosoc_interface_adr;
assign vns_videosoc_interface5_bank_bus_adr = soc_videosoc_videosoc_interface_adr;
assign vns_videosoc_interface6_bank_bus_adr = soc_videosoc_videosoc_interface_adr;
assign vns_videosoc_interface7_bank_bus_adr = soc_videosoc_videosoc_interface_adr;
assign vns_videosoc_interface8_bank_bus_adr = soc_videosoc_videosoc_interface_adr;
assign vns_videosoc_interface9_bank_bus_adr = soc_videosoc_videosoc_interface_adr;
assign vns_videosoc_interface10_bank_bus_adr = soc_videosoc_videosoc_interface_adr;
assign vns_videosoc_interface11_bank_bus_adr = soc_videosoc_videosoc_interface_adr;
assign vns_videosoc_interface12_bank_bus_adr = soc_videosoc_videosoc_interface_adr;
assign vns_videosoc_sram_bus_adr = soc_videosoc_videosoc_interface_adr;
assign vns_videosoc_interface0_bank_bus_we = soc_videosoc_videosoc_interface_we;
assign vns_videosoc_interface1_bank_bus_we = soc_videosoc_videosoc_interface_we;
assign vns_videosoc_interface2_bank_bus_we = soc_videosoc_videosoc_interface_we;
assign vns_videosoc_interface3_bank_bus_we = soc_videosoc_videosoc_interface_we;
assign vns_videosoc_interface4_bank_bus_we = soc_videosoc_videosoc_interface_we;
assign vns_videosoc_interface5_bank_bus_we = soc_videosoc_videosoc_interface_we;
assign vns_videosoc_interface6_bank_bus_we = soc_videosoc_videosoc_interface_we;
assign vns_videosoc_interface7_bank_bus_we = soc_videosoc_videosoc_interface_we;
assign vns_videosoc_interface8_bank_bus_we = soc_videosoc_videosoc_interface_we;
assign vns_videosoc_interface9_bank_bus_we = soc_videosoc_videosoc_interface_we;
assign vns_videosoc_interface10_bank_bus_we = soc_videosoc_videosoc_interface_we;
assign vns_videosoc_interface11_bank_bus_we = soc_videosoc_videosoc_interface_we;
assign vns_videosoc_interface12_bank_bus_we = soc_videosoc_videosoc_interface_we;
assign vns_videosoc_sram_bus_we = soc_videosoc_videosoc_interface_we;
assign vns_videosoc_interface0_bank_bus_dat_w = soc_videosoc_videosoc_interface_dat_w;
assign vns_videosoc_interface1_bank_bus_dat_w = soc_videosoc_videosoc_interface_dat_w;
assign vns_videosoc_interface2_bank_bus_dat_w = soc_videosoc_videosoc_interface_dat_w;
assign vns_videosoc_interface3_bank_bus_dat_w = soc_videosoc_videosoc_interface_dat_w;
assign vns_videosoc_interface4_bank_bus_dat_w = soc_videosoc_videosoc_interface_dat_w;
assign vns_videosoc_interface5_bank_bus_dat_w = soc_videosoc_videosoc_interface_dat_w;
assign vns_videosoc_interface6_bank_bus_dat_w = soc_videosoc_videosoc_interface_dat_w;
assign vns_videosoc_interface7_bank_bus_dat_w = soc_videosoc_videosoc_interface_dat_w;
assign vns_videosoc_interface8_bank_bus_dat_w = soc_videosoc_videosoc_interface_dat_w;
assign vns_videosoc_interface9_bank_bus_dat_w = soc_videosoc_videosoc_interface_dat_w;
assign vns_videosoc_interface10_bank_bus_dat_w = soc_videosoc_videosoc_interface_dat_w;
assign vns_videosoc_interface11_bank_bus_dat_w = soc_videosoc_videosoc_interface_dat_w;
assign vns_videosoc_interface12_bank_bus_dat_w = soc_videosoc_videosoc_interface_dat_w;
assign vns_videosoc_sram_bus_dat_w = soc_videosoc_videosoc_interface_dat_w;
assign soc_videosoc_videosoc_interface_dat_r = (((((((((((((vns_videosoc_interface0_bank_bus_dat_r | vns_videosoc_interface1_bank_bus_dat_r) | vns_videosoc_interface2_bank_bus_dat_r) | vns_videosoc_interface3_bank_bus_dat_r) | vns_videosoc_interface4_bank_bus_dat_r) | vns_videosoc_interface5_bank_bus_dat_r) | vns_videosoc_interface6_bank_bus_dat_r) | vns_videosoc_interface7_bank_bus_dat_r) | vns_videosoc_interface8_bank_bus_dat_r) | vns_videosoc_interface9_bank_bus_dat_r) | vns_videosoc_interface10_bank_bus_dat_r) | vns_videosoc_interface11_bank_bus_dat_r) | vns_videosoc_interface12_bank_bus_dat_r) | vns_videosoc_sram_bus_dat_r);
always @(*) begin
	vns_comb_rhs_array_muxed0 <= 1'd0;
	case (soc_videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed0 <= soc_videosoc_sdram_choose_cmd_valids[0];
		end
		1'd1: begin
			vns_comb_rhs_array_muxed0 <= soc_videosoc_sdram_choose_cmd_valids[1];
		end
		2'd2: begin
			vns_comb_rhs_array_muxed0 <= soc_videosoc_sdram_choose_cmd_valids[2];
		end
		2'd3: begin
			vns_comb_rhs_array_muxed0 <= soc_videosoc_sdram_choose_cmd_valids[3];
		end
		3'd4: begin
			vns_comb_rhs_array_muxed0 <= soc_videosoc_sdram_choose_cmd_valids[4];
		end
		3'd5: begin
			vns_comb_rhs_array_muxed0 <= soc_videosoc_sdram_choose_cmd_valids[5];
		end
		3'd6: begin
			vns_comb_rhs_array_muxed0 <= soc_videosoc_sdram_choose_cmd_valids[6];
		end
		default: begin
			vns_comb_rhs_array_muxed0 <= soc_videosoc_sdram_choose_cmd_valids[7];
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed1 <= 15'd0;
	case (soc_videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed1 <= soc_videosoc_sdram_bankmachine0_cmd_payload_a;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed1 <= soc_videosoc_sdram_bankmachine1_cmd_payload_a;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed1 <= soc_videosoc_sdram_bankmachine2_cmd_payload_a;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed1 <= soc_videosoc_sdram_bankmachine3_cmd_payload_a;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed1 <= soc_videosoc_sdram_bankmachine4_cmd_payload_a;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed1 <= soc_videosoc_sdram_bankmachine5_cmd_payload_a;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed1 <= soc_videosoc_sdram_bankmachine6_cmd_payload_a;
		end
		default: begin
			vns_comb_rhs_array_muxed1 <= soc_videosoc_sdram_bankmachine7_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed2 <= 3'd0;
	case (soc_videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed2 <= soc_videosoc_sdram_bankmachine0_cmd_payload_ba;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed2 <= soc_videosoc_sdram_bankmachine1_cmd_payload_ba;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed2 <= soc_videosoc_sdram_bankmachine2_cmd_payload_ba;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed2 <= soc_videosoc_sdram_bankmachine3_cmd_payload_ba;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed2 <= soc_videosoc_sdram_bankmachine4_cmd_payload_ba;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed2 <= soc_videosoc_sdram_bankmachine5_cmd_payload_ba;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed2 <= soc_videosoc_sdram_bankmachine6_cmd_payload_ba;
		end
		default: begin
			vns_comb_rhs_array_muxed2 <= soc_videosoc_sdram_bankmachine7_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed3 <= 1'd0;
	case (soc_videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed3 <= soc_videosoc_sdram_bankmachine0_cmd_payload_is_read;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed3 <= soc_videosoc_sdram_bankmachine1_cmd_payload_is_read;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed3 <= soc_videosoc_sdram_bankmachine2_cmd_payload_is_read;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed3 <= soc_videosoc_sdram_bankmachine3_cmd_payload_is_read;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed3 <= soc_videosoc_sdram_bankmachine4_cmd_payload_is_read;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed3 <= soc_videosoc_sdram_bankmachine5_cmd_payload_is_read;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed3 <= soc_videosoc_sdram_bankmachine6_cmd_payload_is_read;
		end
		default: begin
			vns_comb_rhs_array_muxed3 <= soc_videosoc_sdram_bankmachine7_cmd_payload_is_read;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed4 <= 1'd0;
	case (soc_videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed4 <= soc_videosoc_sdram_bankmachine0_cmd_payload_is_write;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed4 <= soc_videosoc_sdram_bankmachine1_cmd_payload_is_write;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed4 <= soc_videosoc_sdram_bankmachine2_cmd_payload_is_write;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed4 <= soc_videosoc_sdram_bankmachine3_cmd_payload_is_write;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed4 <= soc_videosoc_sdram_bankmachine4_cmd_payload_is_write;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed4 <= soc_videosoc_sdram_bankmachine5_cmd_payload_is_write;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed4 <= soc_videosoc_sdram_bankmachine6_cmd_payload_is_write;
		end
		default: begin
			vns_comb_rhs_array_muxed4 <= soc_videosoc_sdram_bankmachine7_cmd_payload_is_write;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed5 <= 1'd0;
	case (soc_videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed5 <= soc_videosoc_sdram_bankmachine0_cmd_payload_is_cmd;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed5 <= soc_videosoc_sdram_bankmachine1_cmd_payload_is_cmd;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed5 <= soc_videosoc_sdram_bankmachine2_cmd_payload_is_cmd;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed5 <= soc_videosoc_sdram_bankmachine3_cmd_payload_is_cmd;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed5 <= soc_videosoc_sdram_bankmachine4_cmd_payload_is_cmd;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed5 <= soc_videosoc_sdram_bankmachine5_cmd_payload_is_cmd;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed5 <= soc_videosoc_sdram_bankmachine6_cmd_payload_is_cmd;
		end
		default: begin
			vns_comb_rhs_array_muxed5 <= soc_videosoc_sdram_bankmachine7_cmd_payload_is_cmd;
		end
	endcase
end
always @(*) begin
	vns_comb_t_array_muxed0 <= 1'd0;
	case (soc_videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_t_array_muxed0 <= soc_videosoc_sdram_bankmachine0_cmd_payload_cas;
		end
		1'd1: begin
			vns_comb_t_array_muxed0 <= soc_videosoc_sdram_bankmachine1_cmd_payload_cas;
		end
		2'd2: begin
			vns_comb_t_array_muxed0 <= soc_videosoc_sdram_bankmachine2_cmd_payload_cas;
		end
		2'd3: begin
			vns_comb_t_array_muxed0 <= soc_videosoc_sdram_bankmachine3_cmd_payload_cas;
		end
		3'd4: begin
			vns_comb_t_array_muxed0 <= soc_videosoc_sdram_bankmachine4_cmd_payload_cas;
		end
		3'd5: begin
			vns_comb_t_array_muxed0 <= soc_videosoc_sdram_bankmachine5_cmd_payload_cas;
		end
		3'd6: begin
			vns_comb_t_array_muxed0 <= soc_videosoc_sdram_bankmachine6_cmd_payload_cas;
		end
		default: begin
			vns_comb_t_array_muxed0 <= soc_videosoc_sdram_bankmachine7_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	vns_comb_t_array_muxed1 <= 1'd0;
	case (soc_videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_t_array_muxed1 <= soc_videosoc_sdram_bankmachine0_cmd_payload_ras;
		end
		1'd1: begin
			vns_comb_t_array_muxed1 <= soc_videosoc_sdram_bankmachine1_cmd_payload_ras;
		end
		2'd2: begin
			vns_comb_t_array_muxed1 <= soc_videosoc_sdram_bankmachine2_cmd_payload_ras;
		end
		2'd3: begin
			vns_comb_t_array_muxed1 <= soc_videosoc_sdram_bankmachine3_cmd_payload_ras;
		end
		3'd4: begin
			vns_comb_t_array_muxed1 <= soc_videosoc_sdram_bankmachine4_cmd_payload_ras;
		end
		3'd5: begin
			vns_comb_t_array_muxed1 <= soc_videosoc_sdram_bankmachine5_cmd_payload_ras;
		end
		3'd6: begin
			vns_comb_t_array_muxed1 <= soc_videosoc_sdram_bankmachine6_cmd_payload_ras;
		end
		default: begin
			vns_comb_t_array_muxed1 <= soc_videosoc_sdram_bankmachine7_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	vns_comb_t_array_muxed2 <= 1'd0;
	case (soc_videosoc_sdram_choose_cmd_grant)
		1'd0: begin
			vns_comb_t_array_muxed2 <= soc_videosoc_sdram_bankmachine0_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_t_array_muxed2 <= soc_videosoc_sdram_bankmachine1_cmd_payload_we;
		end
		2'd2: begin
			vns_comb_t_array_muxed2 <= soc_videosoc_sdram_bankmachine2_cmd_payload_we;
		end
		2'd3: begin
			vns_comb_t_array_muxed2 <= soc_videosoc_sdram_bankmachine3_cmd_payload_we;
		end
		3'd4: begin
			vns_comb_t_array_muxed2 <= soc_videosoc_sdram_bankmachine4_cmd_payload_we;
		end
		3'd5: begin
			vns_comb_t_array_muxed2 <= soc_videosoc_sdram_bankmachine5_cmd_payload_we;
		end
		3'd6: begin
			vns_comb_t_array_muxed2 <= soc_videosoc_sdram_bankmachine6_cmd_payload_we;
		end
		default: begin
			vns_comb_t_array_muxed2 <= soc_videosoc_sdram_bankmachine7_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed6 <= 1'd0;
	case (soc_videosoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed6 <= soc_videosoc_sdram_choose_req_valids[0];
		end
		1'd1: begin
			vns_comb_rhs_array_muxed6 <= soc_videosoc_sdram_choose_req_valids[1];
		end
		2'd2: begin
			vns_comb_rhs_array_muxed6 <= soc_videosoc_sdram_choose_req_valids[2];
		end
		2'd3: begin
			vns_comb_rhs_array_muxed6 <= soc_videosoc_sdram_choose_req_valids[3];
		end
		3'd4: begin
			vns_comb_rhs_array_muxed6 <= soc_videosoc_sdram_choose_req_valids[4];
		end
		3'd5: begin
			vns_comb_rhs_array_muxed6 <= soc_videosoc_sdram_choose_req_valids[5];
		end
		3'd6: begin
			vns_comb_rhs_array_muxed6 <= soc_videosoc_sdram_choose_req_valids[6];
		end
		default: begin
			vns_comb_rhs_array_muxed6 <= soc_videosoc_sdram_choose_req_valids[7];
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed7 <= 15'd0;
	case (soc_videosoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed7 <= soc_videosoc_sdram_bankmachine0_cmd_payload_a;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed7 <= soc_videosoc_sdram_bankmachine1_cmd_payload_a;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed7 <= soc_videosoc_sdram_bankmachine2_cmd_payload_a;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed7 <= soc_videosoc_sdram_bankmachine3_cmd_payload_a;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed7 <= soc_videosoc_sdram_bankmachine4_cmd_payload_a;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed7 <= soc_videosoc_sdram_bankmachine5_cmd_payload_a;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed7 <= soc_videosoc_sdram_bankmachine6_cmd_payload_a;
		end
		default: begin
			vns_comb_rhs_array_muxed7 <= soc_videosoc_sdram_bankmachine7_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed8 <= 3'd0;
	case (soc_videosoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed8 <= soc_videosoc_sdram_bankmachine0_cmd_payload_ba;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed8 <= soc_videosoc_sdram_bankmachine1_cmd_payload_ba;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed8 <= soc_videosoc_sdram_bankmachine2_cmd_payload_ba;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed8 <= soc_videosoc_sdram_bankmachine3_cmd_payload_ba;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed8 <= soc_videosoc_sdram_bankmachine4_cmd_payload_ba;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed8 <= soc_videosoc_sdram_bankmachine5_cmd_payload_ba;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed8 <= soc_videosoc_sdram_bankmachine6_cmd_payload_ba;
		end
		default: begin
			vns_comb_rhs_array_muxed8 <= soc_videosoc_sdram_bankmachine7_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed9 <= 1'd0;
	case (soc_videosoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed9 <= soc_videosoc_sdram_bankmachine0_cmd_payload_is_read;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed9 <= soc_videosoc_sdram_bankmachine1_cmd_payload_is_read;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed9 <= soc_videosoc_sdram_bankmachine2_cmd_payload_is_read;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed9 <= soc_videosoc_sdram_bankmachine3_cmd_payload_is_read;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed9 <= soc_videosoc_sdram_bankmachine4_cmd_payload_is_read;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed9 <= soc_videosoc_sdram_bankmachine5_cmd_payload_is_read;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed9 <= soc_videosoc_sdram_bankmachine6_cmd_payload_is_read;
		end
		default: begin
			vns_comb_rhs_array_muxed9 <= soc_videosoc_sdram_bankmachine7_cmd_payload_is_read;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed10 <= 1'd0;
	case (soc_videosoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed10 <= soc_videosoc_sdram_bankmachine0_cmd_payload_is_write;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed10 <= soc_videosoc_sdram_bankmachine1_cmd_payload_is_write;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed10 <= soc_videosoc_sdram_bankmachine2_cmd_payload_is_write;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed10 <= soc_videosoc_sdram_bankmachine3_cmd_payload_is_write;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed10 <= soc_videosoc_sdram_bankmachine4_cmd_payload_is_write;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed10 <= soc_videosoc_sdram_bankmachine5_cmd_payload_is_write;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed10 <= soc_videosoc_sdram_bankmachine6_cmd_payload_is_write;
		end
		default: begin
			vns_comb_rhs_array_muxed10 <= soc_videosoc_sdram_bankmachine7_cmd_payload_is_write;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed11 <= 1'd0;
	case (soc_videosoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed11 <= soc_videosoc_sdram_bankmachine0_cmd_payload_is_cmd;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed11 <= soc_videosoc_sdram_bankmachine1_cmd_payload_is_cmd;
		end
		2'd2: begin
			vns_comb_rhs_array_muxed11 <= soc_videosoc_sdram_bankmachine2_cmd_payload_is_cmd;
		end
		2'd3: begin
			vns_comb_rhs_array_muxed11 <= soc_videosoc_sdram_bankmachine3_cmd_payload_is_cmd;
		end
		3'd4: begin
			vns_comb_rhs_array_muxed11 <= soc_videosoc_sdram_bankmachine4_cmd_payload_is_cmd;
		end
		3'd5: begin
			vns_comb_rhs_array_muxed11 <= soc_videosoc_sdram_bankmachine5_cmd_payload_is_cmd;
		end
		3'd6: begin
			vns_comb_rhs_array_muxed11 <= soc_videosoc_sdram_bankmachine6_cmd_payload_is_cmd;
		end
		default: begin
			vns_comb_rhs_array_muxed11 <= soc_videosoc_sdram_bankmachine7_cmd_payload_is_cmd;
		end
	endcase
end
always @(*) begin
	vns_comb_t_array_muxed3 <= 1'd0;
	case (soc_videosoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_t_array_muxed3 <= soc_videosoc_sdram_bankmachine0_cmd_payload_cas;
		end
		1'd1: begin
			vns_comb_t_array_muxed3 <= soc_videosoc_sdram_bankmachine1_cmd_payload_cas;
		end
		2'd2: begin
			vns_comb_t_array_muxed3 <= soc_videosoc_sdram_bankmachine2_cmd_payload_cas;
		end
		2'd3: begin
			vns_comb_t_array_muxed3 <= soc_videosoc_sdram_bankmachine3_cmd_payload_cas;
		end
		3'd4: begin
			vns_comb_t_array_muxed3 <= soc_videosoc_sdram_bankmachine4_cmd_payload_cas;
		end
		3'd5: begin
			vns_comb_t_array_muxed3 <= soc_videosoc_sdram_bankmachine5_cmd_payload_cas;
		end
		3'd6: begin
			vns_comb_t_array_muxed3 <= soc_videosoc_sdram_bankmachine6_cmd_payload_cas;
		end
		default: begin
			vns_comb_t_array_muxed3 <= soc_videosoc_sdram_bankmachine7_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	vns_comb_t_array_muxed4 <= 1'd0;
	case (soc_videosoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_t_array_muxed4 <= soc_videosoc_sdram_bankmachine0_cmd_payload_ras;
		end
		1'd1: begin
			vns_comb_t_array_muxed4 <= soc_videosoc_sdram_bankmachine1_cmd_payload_ras;
		end
		2'd2: begin
			vns_comb_t_array_muxed4 <= soc_videosoc_sdram_bankmachine2_cmd_payload_ras;
		end
		2'd3: begin
			vns_comb_t_array_muxed4 <= soc_videosoc_sdram_bankmachine3_cmd_payload_ras;
		end
		3'd4: begin
			vns_comb_t_array_muxed4 <= soc_videosoc_sdram_bankmachine4_cmd_payload_ras;
		end
		3'd5: begin
			vns_comb_t_array_muxed4 <= soc_videosoc_sdram_bankmachine5_cmd_payload_ras;
		end
		3'd6: begin
			vns_comb_t_array_muxed4 <= soc_videosoc_sdram_bankmachine6_cmd_payload_ras;
		end
		default: begin
			vns_comb_t_array_muxed4 <= soc_videosoc_sdram_bankmachine7_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	vns_comb_t_array_muxed5 <= 1'd0;
	case (soc_videosoc_sdram_choose_req_grant)
		1'd0: begin
			vns_comb_t_array_muxed5 <= soc_videosoc_sdram_bankmachine0_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_t_array_muxed5 <= soc_videosoc_sdram_bankmachine1_cmd_payload_we;
		end
		2'd2: begin
			vns_comb_t_array_muxed5 <= soc_videosoc_sdram_bankmachine2_cmd_payload_we;
		end
		2'd3: begin
			vns_comb_t_array_muxed5 <= soc_videosoc_sdram_bankmachine3_cmd_payload_we;
		end
		3'd4: begin
			vns_comb_t_array_muxed5 <= soc_videosoc_sdram_bankmachine4_cmd_payload_we;
		end
		3'd5: begin
			vns_comb_t_array_muxed5 <= soc_videosoc_sdram_bankmachine5_cmd_payload_we;
		end
		3'd6: begin
			vns_comb_t_array_muxed5 <= soc_videosoc_sdram_bankmachine6_cmd_payload_we;
		end
		default: begin
			vns_comb_t_array_muxed5 <= soc_videosoc_sdram_bankmachine7_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed12 <= 22'd0;
	case (vns_roundrobin0_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed12 <= vns_rca0;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed12 <= vns_rca1;
		end
		default: begin
			vns_comb_rhs_array_muxed12 <= vns_rca2;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed13 <= 1'd0;
	case (vns_roundrobin0_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed13 <= soc_videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed13 <= soc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed13 <= soc_hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed14 <= 1'd0;
	case (vns_roundrobin0_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed14 <= (((vns_cba0 == 1'd0) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videosoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed14 <= (((vns_cba1 == 1'd0) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed14 <= (((vns_cba2 == 1'd0) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed15 <= 22'd0;
	case (vns_roundrobin1_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed15 <= vns_rca0;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed15 <= vns_rca1;
		end
		default: begin
			vns_comb_rhs_array_muxed15 <= vns_rca2;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed16 <= 1'd0;
	case (vns_roundrobin1_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed16 <= soc_videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed16 <= soc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed16 <= soc_hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed17 <= 1'd0;
	case (vns_roundrobin1_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed17 <= (((vns_cba0 == 1'd1) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videosoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed17 <= (((vns_cba1 == 1'd1) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed17 <= (((vns_cba2 == 1'd1) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed18 <= 22'd0;
	case (vns_roundrobin2_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed18 <= vns_rca0;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed18 <= vns_rca1;
		end
		default: begin
			vns_comb_rhs_array_muxed18 <= vns_rca2;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed19 <= 1'd0;
	case (vns_roundrobin2_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed19 <= soc_videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed19 <= soc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed19 <= soc_hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed20 <= 1'd0;
	case (vns_roundrobin2_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed20 <= (((vns_cba0 == 2'd2) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videosoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed20 <= (((vns_cba1 == 2'd2) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed20 <= (((vns_cba2 == 2'd2) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed21 <= 22'd0;
	case (vns_roundrobin3_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed21 <= vns_rca0;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed21 <= vns_rca1;
		end
		default: begin
			vns_comb_rhs_array_muxed21 <= vns_rca2;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed22 <= 1'd0;
	case (vns_roundrobin3_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed22 <= soc_videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed22 <= soc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed22 <= soc_hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed23 <= 1'd0;
	case (vns_roundrobin3_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed23 <= (((vns_cba0 == 2'd3) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videosoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed23 <= (((vns_cba1 == 2'd3) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed23 <= (((vns_cba2 == 2'd3) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed24 <= 22'd0;
	case (vns_roundrobin4_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed24 <= vns_rca0;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed24 <= vns_rca1;
		end
		default: begin
			vns_comb_rhs_array_muxed24 <= vns_rca2;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed25 <= 1'd0;
	case (vns_roundrobin4_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed25 <= soc_videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed25 <= soc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed25 <= soc_hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed26 <= 1'd0;
	case (vns_roundrobin4_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed26 <= (((vns_cba0 == 3'd4) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videosoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed26 <= (((vns_cba1 == 3'd4) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed26 <= (((vns_cba2 == 3'd4) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed27 <= 22'd0;
	case (vns_roundrobin5_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed27 <= vns_rca0;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed27 <= vns_rca1;
		end
		default: begin
			vns_comb_rhs_array_muxed27 <= vns_rca2;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed28 <= 1'd0;
	case (vns_roundrobin5_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed28 <= soc_videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed28 <= soc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed28 <= soc_hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed29 <= 1'd0;
	case (vns_roundrobin5_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed29 <= (((vns_cba0 == 3'd5) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videosoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed29 <= (((vns_cba1 == 3'd5) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed29 <= (((vns_cba2 == 3'd5) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed30 <= 22'd0;
	case (vns_roundrobin6_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed30 <= vns_rca0;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed30 <= vns_rca1;
		end
		default: begin
			vns_comb_rhs_array_muxed30 <= vns_rca2;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed31 <= 1'd0;
	case (vns_roundrobin6_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed31 <= soc_videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed31 <= soc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed31 <= soc_hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed32 <= 1'd0;
	case (vns_roundrobin6_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed32 <= (((vns_cba0 == 3'd6) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd0))))) & soc_videosoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed32 <= (((vns_cba1 == 3'd6) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed32 <= (((vns_cba2 == 3'd6) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank7_lock & (vns_roundrobin7_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed33 <= 22'd0;
	case (vns_roundrobin7_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed33 <= vns_rca0;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed33 <= vns_rca1;
		end
		default: begin
			vns_comb_rhs_array_muxed33 <= vns_rca2;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed34 <= 1'd0;
	case (vns_roundrobin7_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed34 <= soc_videosoc_port_cmd_payload_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed34 <= soc_litedramcrossbar_cmd_payload_we;
		end
		default: begin
			vns_comb_rhs_array_muxed34 <= soc_hdmi_out0_dram_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed35 <= 1'd0;
	case (vns_roundrobin7_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed35 <= (((vns_cba0 == 3'd7) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd0))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd0))))) & soc_videosoc_port_cmd_valid);
		end
		1'd1: begin
			vns_comb_rhs_array_muxed35 <= (((vns_cba1 == 3'd7) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 1'd1))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 1'd1))))) & soc_litedramcrossbar_cmd_valid);
		end
		default: begin
			vns_comb_rhs_array_muxed35 <= (((vns_cba2 == 3'd7) & (~(((((((1'd0 | (soc_videosoc_sdram_interface_bank0_lock & (vns_roundrobin0_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank1_lock & (vns_roundrobin1_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank2_lock & (vns_roundrobin2_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank3_lock & (vns_roundrobin3_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank4_lock & (vns_roundrobin4_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank5_lock & (vns_roundrobin5_grant == 2'd2))) | (soc_videosoc_sdram_interface_bank6_lock & (vns_roundrobin6_grant == 2'd2))))) & soc_hdmi_out0_dram_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed36 <= 25'd0;
	case (soc_dma_slot_array_current_slot)
		1'd0: begin
			vns_comb_rhs_array_muxed36 <= soc_dma_slot_array_slot0_address;
		end
		default: begin
			vns_comb_rhs_array_muxed36 <= soc_dma_slot_array_slot1_address;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed37 <= 1'd0;
	case (soc_dma_slot_array_current_slot)
		1'd0: begin
			vns_comb_rhs_array_muxed37 <= soc_dma_slot_array_slot0_address_valid;
		end
		default: begin
			vns_comb_rhs_array_muxed37 <= soc_dma_slot_array_slot1_address_valid;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed38 <= 30'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed38 <= soc_videosoc_interface1_wb_sdram_adr;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed39 <= 32'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed39 <= soc_videosoc_interface1_wb_sdram_dat_w;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed40 <= 4'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed40 <= soc_videosoc_interface1_wb_sdram_sel;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed41 <= 1'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed41 <= soc_videosoc_interface1_wb_sdram_cyc;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed42 <= 1'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed42 <= soc_videosoc_interface1_wb_sdram_stb;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed43 <= 1'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed43 <= soc_videosoc_interface1_wb_sdram_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed44 <= 3'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed44 <= soc_videosoc_interface1_wb_sdram_cti;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed45 <= 2'd0;
	case (vns_wb_sdram_con_grant)
		default: begin
			vns_comb_rhs_array_muxed45 <= soc_videosoc_interface1_wb_sdram_bte;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed46 <= 30'd0;
	case (vns_videosoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed46 <= soc_videosoc_videosoc_ibus_adr;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed46 <= soc_videosoc_videosoc_dbus_adr;
		end
		default: begin
			vns_comb_rhs_array_muxed46 <= soc_videosoc_bridge_wishbone_adr;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed47 <= 32'd0;
	case (vns_videosoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed47 <= soc_videosoc_videosoc_ibus_dat_w;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed47 <= soc_videosoc_videosoc_dbus_dat_w;
		end
		default: begin
			vns_comb_rhs_array_muxed47 <= soc_videosoc_bridge_wishbone_dat_w;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed48 <= 4'd0;
	case (vns_videosoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed48 <= soc_videosoc_videosoc_ibus_sel;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed48 <= soc_videosoc_videosoc_dbus_sel;
		end
		default: begin
			vns_comb_rhs_array_muxed48 <= soc_videosoc_bridge_wishbone_sel;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed49 <= 1'd0;
	case (vns_videosoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed49 <= soc_videosoc_videosoc_ibus_cyc;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed49 <= soc_videosoc_videosoc_dbus_cyc;
		end
		default: begin
			vns_comb_rhs_array_muxed49 <= soc_videosoc_bridge_wishbone_cyc;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed50 <= 1'd0;
	case (vns_videosoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed50 <= soc_videosoc_videosoc_ibus_stb;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed50 <= soc_videosoc_videosoc_dbus_stb;
		end
		default: begin
			vns_comb_rhs_array_muxed50 <= soc_videosoc_bridge_wishbone_stb;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed51 <= 1'd0;
	case (vns_videosoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed51 <= soc_videosoc_videosoc_ibus_we;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed51 <= soc_videosoc_videosoc_dbus_we;
		end
		default: begin
			vns_comb_rhs_array_muxed51 <= soc_videosoc_bridge_wishbone_we;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed52 <= 3'd0;
	case (vns_videosoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed52 <= soc_videosoc_videosoc_ibus_cti;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed52 <= soc_videosoc_videosoc_dbus_cti;
		end
		default: begin
			vns_comb_rhs_array_muxed52 <= soc_videosoc_bridge_wishbone_cti;
		end
	endcase
end
always @(*) begin
	vns_comb_rhs_array_muxed53 <= 2'd0;
	case (vns_videosoc_grant)
		1'd0: begin
			vns_comb_rhs_array_muxed53 <= soc_videosoc_videosoc_ibus_bte;
		end
		1'd1: begin
			vns_comb_rhs_array_muxed53 <= soc_videosoc_videosoc_dbus_bte;
		end
		default: begin
			vns_comb_rhs_array_muxed53 <= soc_videosoc_bridge_wishbone_bte;
		end
	endcase
end
always @(*) begin
	vns_sync_f_array_muxed0 <= 10'd0;
	case (soc_hdmi_out0_driver_hdmi_phy_es0_new_c2)
		1'd0: begin
			vns_sync_f_array_muxed0 <= 10'd852;
		end
		1'd1: begin
			vns_sync_f_array_muxed0 <= 8'd171;
		end
		2'd2: begin
			vns_sync_f_array_muxed0 <= 9'd340;
		end
		default: begin
			vns_sync_f_array_muxed0 <= 10'd683;
		end
	endcase
end
always @(*) begin
	vns_sync_f_array_muxed1 <= 10'd0;
	case (soc_hdmi_out0_driver_hdmi_phy_es1_new_c2)
		1'd0: begin
			vns_sync_f_array_muxed1 <= 10'd852;
		end
		1'd1: begin
			vns_sync_f_array_muxed1 <= 8'd171;
		end
		2'd2: begin
			vns_sync_f_array_muxed1 <= 9'd340;
		end
		default: begin
			vns_sync_f_array_muxed1 <= 10'd683;
		end
	endcase
end
always @(*) begin
	vns_sync_f_array_muxed2 <= 10'd0;
	case (soc_hdmi_out0_driver_hdmi_phy_es2_new_c2)
		1'd0: begin
			vns_sync_f_array_muxed2 <= 10'd852;
		end
		1'd1: begin
			vns_sync_f_array_muxed2 <= 8'd171;
		end
		2'd2: begin
			vns_sync_f_array_muxed2 <= 9'd340;
		end
		default: begin
			vns_sync_f_array_muxed2 <= 10'd683;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed0 <= 15'd0;
	case (soc_videosoc_sdram_sel0)
		1'd0: begin
			vns_sync_rhs_array_muxed0 <= soc_videosoc_sdram_nop_a;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed0 <= soc_videosoc_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed0 <= soc_videosoc_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			vns_sync_rhs_array_muxed0 <= soc_videosoc_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed1 <= 3'd0;
	case (soc_videosoc_sdram_sel0)
		1'd0: begin
			vns_sync_rhs_array_muxed1 <= soc_videosoc_sdram_nop_ba;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed1 <= soc_videosoc_sdram_choose_cmd_cmd_payload_ba;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed1 <= soc_videosoc_sdram_choose_req_cmd_payload_ba;
		end
		default: begin
			vns_sync_rhs_array_muxed1 <= soc_videosoc_sdram_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed2 <= 1'd0;
	case (soc_videosoc_sdram_sel0)
		1'd0: begin
			vns_sync_rhs_array_muxed2 <= soc_videosoc_sdram_nop_cas;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed2 <= soc_videosoc_sdram_choose_cmd_cmd_payload_cas;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed2 <= soc_videosoc_sdram_choose_req_cmd_payload_cas;
		end
		default: begin
			vns_sync_rhs_array_muxed2 <= soc_videosoc_sdram_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed3 <= 1'd0;
	case (soc_videosoc_sdram_sel0)
		1'd0: begin
			vns_sync_rhs_array_muxed3 <= soc_videosoc_sdram_nop_ras;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed3 <= soc_videosoc_sdram_choose_cmd_cmd_payload_ras;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed3 <= soc_videosoc_sdram_choose_req_cmd_payload_ras;
		end
		default: begin
			vns_sync_rhs_array_muxed3 <= soc_videosoc_sdram_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed4 <= 1'd0;
	case (soc_videosoc_sdram_sel0)
		1'd0: begin
			vns_sync_rhs_array_muxed4 <= soc_videosoc_sdram_nop_we;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed4 <= soc_videosoc_sdram_choose_cmd_cmd_payload_we;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed4 <= soc_videosoc_sdram_choose_req_cmd_payload_we;
		end
		default: begin
			vns_sync_rhs_array_muxed4 <= soc_videosoc_sdram_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed5 <= 1'd0;
	case (soc_videosoc_sdram_sel0)
		1'd0: begin
			vns_sync_rhs_array_muxed5 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed5 <= (soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed5 <= (soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			vns_sync_rhs_array_muxed5 <= (soc_videosoc_sdram_cmd_valid & soc_videosoc_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed6 <= 1'd0;
	case (soc_videosoc_sdram_sel0)
		1'd0: begin
			vns_sync_rhs_array_muxed6 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed6 <= (soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed6 <= (soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			vns_sync_rhs_array_muxed6 <= (soc_videosoc_sdram_cmd_valid & soc_videosoc_sdram_cmd_payload_is_write);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed7 <= 15'd0;
	case (soc_videosoc_sdram_sel1)
		1'd0: begin
			vns_sync_rhs_array_muxed7 <= soc_videosoc_sdram_nop_a;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed7 <= soc_videosoc_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed7 <= soc_videosoc_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			vns_sync_rhs_array_muxed7 <= soc_videosoc_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed8 <= 3'd0;
	case (soc_videosoc_sdram_sel1)
		1'd0: begin
			vns_sync_rhs_array_muxed8 <= soc_videosoc_sdram_nop_ba;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed8 <= soc_videosoc_sdram_choose_cmd_cmd_payload_ba;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed8 <= soc_videosoc_sdram_choose_req_cmd_payload_ba;
		end
		default: begin
			vns_sync_rhs_array_muxed8 <= soc_videosoc_sdram_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed9 <= 1'd0;
	case (soc_videosoc_sdram_sel1)
		1'd0: begin
			vns_sync_rhs_array_muxed9 <= soc_videosoc_sdram_nop_cas;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed9 <= soc_videosoc_sdram_choose_cmd_cmd_payload_cas;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed9 <= soc_videosoc_sdram_choose_req_cmd_payload_cas;
		end
		default: begin
			vns_sync_rhs_array_muxed9 <= soc_videosoc_sdram_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed10 <= 1'd0;
	case (soc_videosoc_sdram_sel1)
		1'd0: begin
			vns_sync_rhs_array_muxed10 <= soc_videosoc_sdram_nop_ras;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed10 <= soc_videosoc_sdram_choose_cmd_cmd_payload_ras;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed10 <= soc_videosoc_sdram_choose_req_cmd_payload_ras;
		end
		default: begin
			vns_sync_rhs_array_muxed10 <= soc_videosoc_sdram_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed11 <= 1'd0;
	case (soc_videosoc_sdram_sel1)
		1'd0: begin
			vns_sync_rhs_array_muxed11 <= soc_videosoc_sdram_nop_we;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed11 <= soc_videosoc_sdram_choose_cmd_cmd_payload_we;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed11 <= soc_videosoc_sdram_choose_req_cmd_payload_we;
		end
		default: begin
			vns_sync_rhs_array_muxed11 <= soc_videosoc_sdram_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed12 <= 1'd0;
	case (soc_videosoc_sdram_sel1)
		1'd0: begin
			vns_sync_rhs_array_muxed12 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed12 <= (soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed12 <= (soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			vns_sync_rhs_array_muxed12 <= (soc_videosoc_sdram_cmd_valid & soc_videosoc_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed13 <= 1'd0;
	case (soc_videosoc_sdram_sel1)
		1'd0: begin
			vns_sync_rhs_array_muxed13 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed13 <= (soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed13 <= (soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			vns_sync_rhs_array_muxed13 <= (soc_videosoc_sdram_cmd_valid & soc_videosoc_sdram_cmd_payload_is_write);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed14 <= 15'd0;
	case (soc_videosoc_sdram_sel2)
		1'd0: begin
			vns_sync_rhs_array_muxed14 <= soc_videosoc_sdram_nop_a;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed14 <= soc_videosoc_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed14 <= soc_videosoc_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			vns_sync_rhs_array_muxed14 <= soc_videosoc_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed15 <= 3'd0;
	case (soc_videosoc_sdram_sel2)
		1'd0: begin
			vns_sync_rhs_array_muxed15 <= soc_videosoc_sdram_nop_ba;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed15 <= soc_videosoc_sdram_choose_cmd_cmd_payload_ba;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed15 <= soc_videosoc_sdram_choose_req_cmd_payload_ba;
		end
		default: begin
			vns_sync_rhs_array_muxed15 <= soc_videosoc_sdram_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed16 <= 1'd0;
	case (soc_videosoc_sdram_sel2)
		1'd0: begin
			vns_sync_rhs_array_muxed16 <= soc_videosoc_sdram_nop_cas;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed16 <= soc_videosoc_sdram_choose_cmd_cmd_payload_cas;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed16 <= soc_videosoc_sdram_choose_req_cmd_payload_cas;
		end
		default: begin
			vns_sync_rhs_array_muxed16 <= soc_videosoc_sdram_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed17 <= 1'd0;
	case (soc_videosoc_sdram_sel2)
		1'd0: begin
			vns_sync_rhs_array_muxed17 <= soc_videosoc_sdram_nop_ras;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed17 <= soc_videosoc_sdram_choose_cmd_cmd_payload_ras;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed17 <= soc_videosoc_sdram_choose_req_cmd_payload_ras;
		end
		default: begin
			vns_sync_rhs_array_muxed17 <= soc_videosoc_sdram_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed18 <= 1'd0;
	case (soc_videosoc_sdram_sel2)
		1'd0: begin
			vns_sync_rhs_array_muxed18 <= soc_videosoc_sdram_nop_we;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed18 <= soc_videosoc_sdram_choose_cmd_cmd_payload_we;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed18 <= soc_videosoc_sdram_choose_req_cmd_payload_we;
		end
		default: begin
			vns_sync_rhs_array_muxed18 <= soc_videosoc_sdram_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed19 <= 1'd0;
	case (soc_videosoc_sdram_sel2)
		1'd0: begin
			vns_sync_rhs_array_muxed19 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed19 <= (soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed19 <= (soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			vns_sync_rhs_array_muxed19 <= (soc_videosoc_sdram_cmd_valid & soc_videosoc_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed20 <= 1'd0;
	case (soc_videosoc_sdram_sel2)
		1'd0: begin
			vns_sync_rhs_array_muxed20 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed20 <= (soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed20 <= (soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			vns_sync_rhs_array_muxed20 <= (soc_videosoc_sdram_cmd_valid & soc_videosoc_sdram_cmd_payload_is_write);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed21 <= 15'd0;
	case (soc_videosoc_sdram_sel3)
		1'd0: begin
			vns_sync_rhs_array_muxed21 <= soc_videosoc_sdram_nop_a;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed21 <= soc_videosoc_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed21 <= soc_videosoc_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			vns_sync_rhs_array_muxed21 <= soc_videosoc_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed22 <= 3'd0;
	case (soc_videosoc_sdram_sel3)
		1'd0: begin
			vns_sync_rhs_array_muxed22 <= soc_videosoc_sdram_nop_ba;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed22 <= soc_videosoc_sdram_choose_cmd_cmd_payload_ba;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed22 <= soc_videosoc_sdram_choose_req_cmd_payload_ba;
		end
		default: begin
			vns_sync_rhs_array_muxed22 <= soc_videosoc_sdram_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed23 <= 1'd0;
	case (soc_videosoc_sdram_sel3)
		1'd0: begin
			vns_sync_rhs_array_muxed23 <= soc_videosoc_sdram_nop_cas;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed23 <= soc_videosoc_sdram_choose_cmd_cmd_payload_cas;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed23 <= soc_videosoc_sdram_choose_req_cmd_payload_cas;
		end
		default: begin
			vns_sync_rhs_array_muxed23 <= soc_videosoc_sdram_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed24 <= 1'd0;
	case (soc_videosoc_sdram_sel3)
		1'd0: begin
			vns_sync_rhs_array_muxed24 <= soc_videosoc_sdram_nop_ras;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed24 <= soc_videosoc_sdram_choose_cmd_cmd_payload_ras;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed24 <= soc_videosoc_sdram_choose_req_cmd_payload_ras;
		end
		default: begin
			vns_sync_rhs_array_muxed24 <= soc_videosoc_sdram_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed25 <= 1'd0;
	case (soc_videosoc_sdram_sel3)
		1'd0: begin
			vns_sync_rhs_array_muxed25 <= soc_videosoc_sdram_nop_we;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed25 <= soc_videosoc_sdram_choose_cmd_cmd_payload_we;
		end
		2'd2: begin
			vns_sync_rhs_array_muxed25 <= soc_videosoc_sdram_choose_req_cmd_payload_we;
		end
		default: begin
			vns_sync_rhs_array_muxed25 <= soc_videosoc_sdram_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed26 <= 1'd0;
	case (soc_videosoc_sdram_sel3)
		1'd0: begin
			vns_sync_rhs_array_muxed26 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed26 <= (soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed26 <= (soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			vns_sync_rhs_array_muxed26 <= (soc_videosoc_sdram_cmd_valid & soc_videosoc_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	vns_sync_rhs_array_muxed27 <= 1'd0;
	case (soc_videosoc_sdram_sel3)
		1'd0: begin
			vns_sync_rhs_array_muxed27 <= 1'd0;
		end
		1'd1: begin
			vns_sync_rhs_array_muxed27 <= (soc_videosoc_sdram_choose_cmd_cmd_valid & soc_videosoc_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			vns_sync_rhs_array_muxed27 <= (soc_videosoc_sdram_choose_req_cmd_valid & soc_videosoc_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			vns_sync_rhs_array_muxed27 <= (soc_videosoc_sdram_cmd_valid & soc_videosoc_sdram_cmd_payload_is_write);
		end
	endcase
end
assign vns_xilinxasyncresetsynchronizerimpl0 = ((~soc_videosoc_pll_locked) | (~cpu_reset));
assign vns_xilinxasyncresetsynchronizerimpl1 = ((~soc_videosoc_pll_locked) | (~cpu_reset));
assign vns_xilinxasyncresetsynchronizerimpl2 = ((~soc_videosoc_pll_locked) | (~cpu_reset));
assign soc_videosoc_uart_phy_rx = vns_xilinxmultiregimpl0_regs1;
assign soc_ethphy_status = vns_xilinxmultiregimpl1_regs1;
assign soc_ethmac_tx_cdc_produce_rdomain = vns_xilinxmultiregimpl2_regs1;
assign soc_ethmac_tx_cdc_consume_wdomain = vns_xilinxmultiregimpl3_regs1;
assign soc_ethmac_rx_cdc_produce_rdomain = vns_xilinxmultiregimpl4_regs1;
assign soc_ethmac_rx_cdc_consume_wdomain = vns_xilinxmultiregimpl5_regs1;
assign soc_edid_scl_raw = vns_xilinxmultiregimpl6_regs1;
assign soc_edid_sda_raw = vns_xilinxmultiregimpl7_regs1;
assign soc_locked = vns_xilinxmultiregimpl8_regs1;
assign vns_xilinxasyncresetsynchronizerimpl5 = (~soc_mmcm_locked);
assign vns_xilinxasyncresetsynchronizerimpl6 = (~soc_mmcm_locked);
assign soc_s7datacapture0_do_delay_rst_toggle_o = vns_xilinxmultiregimpl9_regs1;
assign soc_s7datacapture0_do_delay_master_inc_toggle_o = vns_xilinxmultiregimpl10_regs1;
assign soc_s7datacapture0_do_delay_master_dec_toggle_o = vns_xilinxmultiregimpl11_regs1;
assign soc_s7datacapture0_do_delay_slave_inc_toggle_o = vns_xilinxmultiregimpl12_regs1;
assign soc_s7datacapture0_do_delay_slave_dec_toggle_o = vns_xilinxmultiregimpl13_regs1;
assign soc_s7datacapture0_status = vns_xilinxmultiregimpl14_regs1;
assign soc_s7datacapture0_do_reset_lateness_toggle_o = vns_xilinxmultiregimpl15_regs1;
assign soc_charsync0_char_synced_status = vns_xilinxmultiregimpl16_regs1;
assign soc_charsync0_ctl_pos_status = vns_xilinxmultiregimpl17_regs1;
assign soc_wer0_toggle_o = vns_xilinxmultiregimpl18_regs1;
assign soc_s7datacapture1_do_delay_rst_toggle_o = vns_xilinxmultiregimpl19_regs1;
assign soc_s7datacapture1_do_delay_master_inc_toggle_o = vns_xilinxmultiregimpl20_regs1;
assign soc_s7datacapture1_do_delay_master_dec_toggle_o = vns_xilinxmultiregimpl21_regs1;
assign soc_s7datacapture1_do_delay_slave_inc_toggle_o = vns_xilinxmultiregimpl22_regs1;
assign soc_s7datacapture1_do_delay_slave_dec_toggle_o = vns_xilinxmultiregimpl23_regs1;
assign soc_s7datacapture1_status = vns_xilinxmultiregimpl24_regs1;
assign soc_s7datacapture1_do_reset_lateness_toggle_o = vns_xilinxmultiregimpl25_regs1;
assign soc_charsync1_char_synced_status = vns_xilinxmultiregimpl26_regs1;
assign soc_charsync1_ctl_pos_status = vns_xilinxmultiregimpl27_regs1;
assign soc_wer1_toggle_o = vns_xilinxmultiregimpl28_regs1;
assign soc_s7datacapture2_do_delay_rst_toggle_o = vns_xilinxmultiregimpl29_regs1;
assign soc_s7datacapture2_do_delay_master_inc_toggle_o = vns_xilinxmultiregimpl30_regs1;
assign soc_s7datacapture2_do_delay_master_dec_toggle_o = vns_xilinxmultiregimpl31_regs1;
assign soc_s7datacapture2_do_delay_slave_inc_toggle_o = vns_xilinxmultiregimpl32_regs1;
assign soc_s7datacapture2_do_delay_slave_dec_toggle_o = vns_xilinxmultiregimpl33_regs1;
assign soc_s7datacapture2_status = vns_xilinxmultiregimpl34_regs1;
assign soc_s7datacapture2_do_reset_lateness_toggle_o = vns_xilinxmultiregimpl35_regs1;
assign soc_charsync2_char_synced_status = vns_xilinxmultiregimpl36_regs1;
assign soc_charsync2_ctl_pos_status = vns_xilinxmultiregimpl37_regs1;
assign soc_wer2_toggle_o = vns_xilinxmultiregimpl38_regs1;
assign soc_chansync_status = vns_xilinxmultiregimpl39_regs1;
assign soc_resdetection_hres_status = vns_xilinxmultiregimpl40_regs1;
assign soc_resdetection_vres_status = vns_xilinxmultiregimpl41_regs1;
assign soc_frame_fifo_produce_rdomain = vns_xilinxmultiregimpl42_regs1;
assign soc_frame_fifo_consume_wdomain = vns_xilinxmultiregimpl43_regs1;
assign soc_frame_sys_overflow = vns_xilinxmultiregimpl44_regs1;
assign soc_frame_overflow_reset_toggle_o = vns_xilinxmultiregimpl45_regs1;
assign soc_frame_overflow_reset_ack_toggle_o = vns_xilinxmultiregimpl46_regs1;
assign soc_hdmi_in0_freq_gray_decoder_i = vns_xilinxmultiregimpl47_regs1;
assign soc_hdmi_out0_dram_port_cmd_fifo_produce_rdomain = vns_xilinxmultiregimpl48_regs1;
assign soc_hdmi_out0_dram_port_cmd_fifo_consume_wdomain = vns_xilinxmultiregimpl49_regs1;
assign soc_hdmi_out0_dram_port_rdata_fifo_produce_rdomain = vns_xilinxmultiregimpl50_regs1;
assign soc_hdmi_out0_dram_port_rdata_fifo_consume_wdomain = vns_xilinxmultiregimpl51_regs1;
assign soc_hdmi_out0_core_initiator_cdc_produce_rdomain = vns_xilinxmultiregimpl52_regs1;
assign soc_hdmi_out0_core_initiator_cdc_consume_wdomain = vns_xilinxmultiregimpl53_regs1;
assign soc_hdmi_out0_core_underflow_enable = vns_xilinxmultiregimpl54_regs1;
assign soc_hdmi_out0_core_toggle_o = vns_xilinxmultiregimpl55_regs1;

always @(posedge clk200_clk) begin
	if ((soc_videosoc_reset_counter != 1'd0)) begin
		soc_videosoc_reset_counter <= (soc_videosoc_reset_counter - 1'd1);
	end else begin
		soc_videosoc_ic_reset <= 1'd0;
	end
	if (clk200_rst) begin
		soc_videosoc_reset_counter <= 4'd15;
		soc_videosoc_ic_reset <= 1'd1;
	end
end

always @(posedge data0_cap_read_clk) begin
	if ((soc_s7datacapture0_gearbox_rdpointer == 3'd7)) begin
		soc_s7datacapture0_gearbox_rdpointer <= 1'd0;
	end else begin
		soc_s7datacapture0_gearbox_rdpointer <= (soc_s7datacapture0_gearbox_rdpointer + 1'd1);
	end
	case (soc_s7datacapture0_gearbox_rdpointer)
		1'd0: begin
			soc_s7datacapture0_gearbox_o <= soc_s7datacapture0_gearbox_storage[9:0];
		end
		1'd1: begin
			soc_s7datacapture0_gearbox_o <= soc_s7datacapture0_gearbox_storage[19:10];
		end
		2'd2: begin
			soc_s7datacapture0_gearbox_o <= soc_s7datacapture0_gearbox_storage[29:20];
		end
		2'd3: begin
			soc_s7datacapture0_gearbox_o <= soc_s7datacapture0_gearbox_storage[39:30];
		end
		3'd4: begin
			soc_s7datacapture0_gearbox_o <= soc_s7datacapture0_gearbox_storage[49:40];
		end
		3'd5: begin
			soc_s7datacapture0_gearbox_o <= soc_s7datacapture0_gearbox_storage[59:50];
		end
		3'd6: begin
			soc_s7datacapture0_gearbox_o <= soc_s7datacapture0_gearbox_storage[69:60];
		end
		3'd7: begin
			soc_s7datacapture0_gearbox_o <= soc_s7datacapture0_gearbox_storage[79:70];
		end
	endcase
	if (data0_cap_read_rst) begin
		soc_s7datacapture0_gearbox_rdpointer <= 3'd0;
	end
end

always @(posedge data0_cap_write_clk) begin
	if ((soc_s7datacapture0_gearbox_wrpointer == 4'd9)) begin
		soc_s7datacapture0_gearbox_wrpointer <= 1'd0;
	end else begin
		soc_s7datacapture0_gearbox_wrpointer <= (soc_s7datacapture0_gearbox_wrpointer + 1'd1);
	end
	case (soc_s7datacapture0_gearbox_wrpointer)
		1'd0: begin
			soc_s7datacapture0_gearbox_storage[7:0] <= soc_s7datacapture0_gearbox_i;
		end
		1'd1: begin
			soc_s7datacapture0_gearbox_storage[15:8] <= soc_s7datacapture0_gearbox_i;
		end
		2'd2: begin
			soc_s7datacapture0_gearbox_storage[23:16] <= soc_s7datacapture0_gearbox_i;
		end
		2'd3: begin
			soc_s7datacapture0_gearbox_storage[31:24] <= soc_s7datacapture0_gearbox_i;
		end
		3'd4: begin
			soc_s7datacapture0_gearbox_storage[39:32] <= soc_s7datacapture0_gearbox_i;
		end
		3'd5: begin
			soc_s7datacapture0_gearbox_storage[47:40] <= soc_s7datacapture0_gearbox_i;
		end
		3'd6: begin
			soc_s7datacapture0_gearbox_storage[55:48] <= soc_s7datacapture0_gearbox_i;
		end
		3'd7: begin
			soc_s7datacapture0_gearbox_storage[63:56] <= soc_s7datacapture0_gearbox_i;
		end
		4'd8: begin
			soc_s7datacapture0_gearbox_storage[71:64] <= soc_s7datacapture0_gearbox_i;
		end
		4'd9: begin
			soc_s7datacapture0_gearbox_storage[79:72] <= soc_s7datacapture0_gearbox_i;
		end
	endcase
	if (data0_cap_write_rst) begin
		soc_s7datacapture0_gearbox_wrpointer <= 4'd5;
	end
end

always @(posedge data1_cap_read_clk) begin
	if ((soc_s7datacapture1_gearbox_rdpointer == 3'd7)) begin
		soc_s7datacapture1_gearbox_rdpointer <= 1'd0;
	end else begin
		soc_s7datacapture1_gearbox_rdpointer <= (soc_s7datacapture1_gearbox_rdpointer + 1'd1);
	end
	case (soc_s7datacapture1_gearbox_rdpointer)
		1'd0: begin
			soc_s7datacapture1_gearbox_o <= soc_s7datacapture1_gearbox_storage[9:0];
		end
		1'd1: begin
			soc_s7datacapture1_gearbox_o <= soc_s7datacapture1_gearbox_storage[19:10];
		end
		2'd2: begin
			soc_s7datacapture1_gearbox_o <= soc_s7datacapture1_gearbox_storage[29:20];
		end
		2'd3: begin
			soc_s7datacapture1_gearbox_o <= soc_s7datacapture1_gearbox_storage[39:30];
		end
		3'd4: begin
			soc_s7datacapture1_gearbox_o <= soc_s7datacapture1_gearbox_storage[49:40];
		end
		3'd5: begin
			soc_s7datacapture1_gearbox_o <= soc_s7datacapture1_gearbox_storage[59:50];
		end
		3'd6: begin
			soc_s7datacapture1_gearbox_o <= soc_s7datacapture1_gearbox_storage[69:60];
		end
		3'd7: begin
			soc_s7datacapture1_gearbox_o <= soc_s7datacapture1_gearbox_storage[79:70];
		end
	endcase
	if (data1_cap_read_rst) begin
		soc_s7datacapture1_gearbox_rdpointer <= 3'd0;
	end
end

always @(posedge data1_cap_write_clk) begin
	if ((soc_s7datacapture1_gearbox_wrpointer == 4'd9)) begin
		soc_s7datacapture1_gearbox_wrpointer <= 1'd0;
	end else begin
		soc_s7datacapture1_gearbox_wrpointer <= (soc_s7datacapture1_gearbox_wrpointer + 1'd1);
	end
	case (soc_s7datacapture1_gearbox_wrpointer)
		1'd0: begin
			soc_s7datacapture1_gearbox_storage[7:0] <= soc_s7datacapture1_gearbox_i;
		end
		1'd1: begin
			soc_s7datacapture1_gearbox_storage[15:8] <= soc_s7datacapture1_gearbox_i;
		end
		2'd2: begin
			soc_s7datacapture1_gearbox_storage[23:16] <= soc_s7datacapture1_gearbox_i;
		end
		2'd3: begin
			soc_s7datacapture1_gearbox_storage[31:24] <= soc_s7datacapture1_gearbox_i;
		end
		3'd4: begin
			soc_s7datacapture1_gearbox_storage[39:32] <= soc_s7datacapture1_gearbox_i;
		end
		3'd5: begin
			soc_s7datacapture1_gearbox_storage[47:40] <= soc_s7datacapture1_gearbox_i;
		end
		3'd6: begin
			soc_s7datacapture1_gearbox_storage[55:48] <= soc_s7datacapture1_gearbox_i;
		end
		3'd7: begin
			soc_s7datacapture1_gearbox_storage[63:56] <= soc_s7datacapture1_gearbox_i;
		end
		4'd8: begin
			soc_s7datacapture1_gearbox_storage[71:64] <= soc_s7datacapture1_gearbox_i;
		end
		4'd9: begin
			soc_s7datacapture1_gearbox_storage[79:72] <= soc_s7datacapture1_gearbox_i;
		end
	endcase
	if (data1_cap_write_rst) begin
		soc_s7datacapture1_gearbox_wrpointer <= 4'd5;
	end
end

always @(posedge data2_cap_read_clk) begin
	if ((soc_s7datacapture2_gearbox_rdpointer == 3'd7)) begin
		soc_s7datacapture2_gearbox_rdpointer <= 1'd0;
	end else begin
		soc_s7datacapture2_gearbox_rdpointer <= (soc_s7datacapture2_gearbox_rdpointer + 1'd1);
	end
	case (soc_s7datacapture2_gearbox_rdpointer)
		1'd0: begin
			soc_s7datacapture2_gearbox_o <= soc_s7datacapture2_gearbox_storage[9:0];
		end
		1'd1: begin
			soc_s7datacapture2_gearbox_o <= soc_s7datacapture2_gearbox_storage[19:10];
		end
		2'd2: begin
			soc_s7datacapture2_gearbox_o <= soc_s7datacapture2_gearbox_storage[29:20];
		end
		2'd3: begin
			soc_s7datacapture2_gearbox_o <= soc_s7datacapture2_gearbox_storage[39:30];
		end
		3'd4: begin
			soc_s7datacapture2_gearbox_o <= soc_s7datacapture2_gearbox_storage[49:40];
		end
		3'd5: begin
			soc_s7datacapture2_gearbox_o <= soc_s7datacapture2_gearbox_storage[59:50];
		end
		3'd6: begin
			soc_s7datacapture2_gearbox_o <= soc_s7datacapture2_gearbox_storage[69:60];
		end
		3'd7: begin
			soc_s7datacapture2_gearbox_o <= soc_s7datacapture2_gearbox_storage[79:70];
		end
	endcase
	if (data2_cap_read_rst) begin
		soc_s7datacapture2_gearbox_rdpointer <= 3'd0;
	end
end

always @(posedge data2_cap_write_clk) begin
	if ((soc_s7datacapture2_gearbox_wrpointer == 4'd9)) begin
		soc_s7datacapture2_gearbox_wrpointer <= 1'd0;
	end else begin
		soc_s7datacapture2_gearbox_wrpointer <= (soc_s7datacapture2_gearbox_wrpointer + 1'd1);
	end
	case (soc_s7datacapture2_gearbox_wrpointer)
		1'd0: begin
			soc_s7datacapture2_gearbox_storage[7:0] <= soc_s7datacapture2_gearbox_i;
		end
		1'd1: begin
			soc_s7datacapture2_gearbox_storage[15:8] <= soc_s7datacapture2_gearbox_i;
		end
		2'd2: begin
			soc_s7datacapture2_gearbox_storage[23:16] <= soc_s7datacapture2_gearbox_i;
		end
		2'd3: begin
			soc_s7datacapture2_gearbox_storage[31:24] <= soc_s7datacapture2_gearbox_i;
		end
		3'd4: begin
			soc_s7datacapture2_gearbox_storage[39:32] <= soc_s7datacapture2_gearbox_i;
		end
		3'd5: begin
			soc_s7datacapture2_gearbox_storage[47:40] <= soc_s7datacapture2_gearbox_i;
		end
		3'd6: begin
			soc_s7datacapture2_gearbox_storage[55:48] <= soc_s7datacapture2_gearbox_i;
		end
		3'd7: begin
			soc_s7datacapture2_gearbox_storage[63:56] <= soc_s7datacapture2_gearbox_i;
		end
		4'd8: begin
			soc_s7datacapture2_gearbox_storage[71:64] <= soc_s7datacapture2_gearbox_i;
		end
		4'd9: begin
			soc_s7datacapture2_gearbox_storage[79:72] <= soc_s7datacapture2_gearbox_i;
		end
	endcase
	if (data2_cap_write_rst) begin
		soc_s7datacapture2_gearbox_wrpointer <= 4'd5;
	end
end

always @(posedge eth_rx_clk) begin
	soc_ethphy_rx_ctl_d <= soc_ethphy_rx_ctl;
	soc_ethphy_source_valid <= soc_ethphy_rx_ctl;
	soc_ethphy_source_payload_data <= soc_ethphy_rx_data;
	if (soc_ethmac_rx_gap_checker_counter_reset) begin
		soc_ethmac_rx_gap_checker_counter <= 1'd0;
	end else begin
		if (soc_ethmac_rx_gap_checker_counter_ce) begin
			soc_ethmac_rx_gap_checker_counter <= (soc_ethmac_rx_gap_checker_counter + 1'd1);
		end
	end
	vns_clockdomainsrenamer1_state <= vns_clockdomainsrenamer1_next_state;
	if (soc_ethmac_preamble_checker_clr_cnt) begin
		soc_ethmac_preamble_checker_cnt <= 1'd0;
	end else begin
		if (soc_ethmac_preamble_checker_inc_cnt) begin
			soc_ethmac_preamble_checker_cnt <= (soc_ethmac_preamble_checker_cnt + 1'd1);
		end
	end
	if (soc_ethmac_preamble_checker_clr_discard) begin
		soc_ethmac_preamble_checker_discard <= 1'd0;
	end else begin
		if (soc_ethmac_preamble_checker_set_discard) begin
			soc_ethmac_preamble_checker_discard <= 1'd1;
		end
	end
	vns_clockdomainsrenamer3_state <= vns_clockdomainsrenamer3_next_state;
	if (soc_ethmac_crc32_checker_crc_ce) begin
		soc_ethmac_crc32_checker_crc_reg <= soc_ethmac_crc32_checker_crc_next;
	end
	if (soc_ethmac_crc32_checker_crc_reset) begin
		soc_ethmac_crc32_checker_crc_reg <= 32'd4294967295;
	end
	if (((soc_ethmac_crc32_checker_syncfifo_syncfifo_we & soc_ethmac_crc32_checker_syncfifo_syncfifo_writable) & (~soc_ethmac_crc32_checker_syncfifo_replace))) begin
		if ((soc_ethmac_crc32_checker_syncfifo_produce == 3'd4)) begin
			soc_ethmac_crc32_checker_syncfifo_produce <= 1'd0;
		end else begin
			soc_ethmac_crc32_checker_syncfifo_produce <= (soc_ethmac_crc32_checker_syncfifo_produce + 1'd1);
		end
	end
	if (soc_ethmac_crc32_checker_syncfifo_do_read) begin
		if ((soc_ethmac_crc32_checker_syncfifo_consume == 3'd4)) begin
			soc_ethmac_crc32_checker_syncfifo_consume <= 1'd0;
		end else begin
			soc_ethmac_crc32_checker_syncfifo_consume <= (soc_ethmac_crc32_checker_syncfifo_consume + 1'd1);
		end
	end
	if (((soc_ethmac_crc32_checker_syncfifo_syncfifo_we & soc_ethmac_crc32_checker_syncfifo_syncfifo_writable) & (~soc_ethmac_crc32_checker_syncfifo_replace))) begin
		if ((~soc_ethmac_crc32_checker_syncfifo_do_read)) begin
			soc_ethmac_crc32_checker_syncfifo_level <= (soc_ethmac_crc32_checker_syncfifo_level + 1'd1);
		end
	end else begin
		if (soc_ethmac_crc32_checker_syncfifo_do_read) begin
			soc_ethmac_crc32_checker_syncfifo_level <= (soc_ethmac_crc32_checker_syncfifo_level - 1'd1);
		end
	end
	if (soc_ethmac_crc32_checker_fifo_reset) begin
		soc_ethmac_crc32_checker_syncfifo_level <= 3'd0;
		soc_ethmac_crc32_checker_syncfifo_produce <= 3'd0;
		soc_ethmac_crc32_checker_syncfifo_consume <= 3'd0;
	end
	vns_clockdomainsrenamer5_state <= vns_clockdomainsrenamer5_next_state;
	if (soc_ethmac_rx_converter_converter_source_ready) begin
		soc_ethmac_rx_converter_converter_strobe_all <= 1'd0;
	end
	if (soc_ethmac_rx_converter_converter_load_part) begin
		if (((soc_ethmac_rx_converter_converter_demux == 2'd3) | soc_ethmac_rx_converter_converter_sink_last)) begin
			soc_ethmac_rx_converter_converter_demux <= 1'd0;
			soc_ethmac_rx_converter_converter_strobe_all <= 1'd1;
		end else begin
			soc_ethmac_rx_converter_converter_demux <= (soc_ethmac_rx_converter_converter_demux + 1'd1);
		end
	end
	if ((soc_ethmac_rx_converter_converter_source_valid & soc_ethmac_rx_converter_converter_source_ready)) begin
		if ((soc_ethmac_rx_converter_converter_sink_valid & soc_ethmac_rx_converter_converter_sink_ready)) begin
			soc_ethmac_rx_converter_converter_source_first <= soc_ethmac_rx_converter_converter_sink_first;
			soc_ethmac_rx_converter_converter_source_last <= soc_ethmac_rx_converter_converter_sink_last;
		end else begin
			soc_ethmac_rx_converter_converter_source_first <= 1'd0;
			soc_ethmac_rx_converter_converter_source_last <= 1'd0;
		end
	end else begin
		if ((soc_ethmac_rx_converter_converter_sink_valid & soc_ethmac_rx_converter_converter_sink_ready)) begin
			soc_ethmac_rx_converter_converter_source_first <= (soc_ethmac_rx_converter_converter_sink_first | soc_ethmac_rx_converter_converter_source_first);
			soc_ethmac_rx_converter_converter_source_last <= (soc_ethmac_rx_converter_converter_sink_last | soc_ethmac_rx_converter_converter_source_last);
		end
	end
	if (soc_ethmac_rx_converter_converter_load_part) begin
		case (soc_ethmac_rx_converter_converter_demux)
			1'd0: begin
				soc_ethmac_rx_converter_converter_source_payload_data[39:30] <= soc_ethmac_rx_converter_converter_sink_payload_data;
			end
			1'd1: begin
				soc_ethmac_rx_converter_converter_source_payload_data[29:20] <= soc_ethmac_rx_converter_converter_sink_payload_data;
			end
			2'd2: begin
				soc_ethmac_rx_converter_converter_source_payload_data[19:10] <= soc_ethmac_rx_converter_converter_sink_payload_data;
			end
			2'd3: begin
				soc_ethmac_rx_converter_converter_source_payload_data[9:0] <= soc_ethmac_rx_converter_converter_sink_payload_data;
			end
		endcase
	end
	if (soc_ethmac_rx_converter_converter_load_part) begin
		soc_ethmac_rx_converter_converter_source_payload_valid_token_count <= (soc_ethmac_rx_converter_converter_demux + 1'd1);
	end
	soc_ethmac_rx_cdc_graycounter0_q_binary <= soc_ethmac_rx_cdc_graycounter0_q_next_binary;
	soc_ethmac_rx_cdc_graycounter0_q <= soc_ethmac_rx_cdc_graycounter0_q_next;
	if (eth_rx_rst) begin
		soc_ethphy_source_valid <= 1'd0;
		soc_ethphy_rx_ctl_d <= 1'd0;
		soc_ethmac_crc32_checker_crc_reg <= 32'd4294967295;
		soc_ethmac_crc32_checker_syncfifo_level <= 3'd0;
		soc_ethmac_crc32_checker_syncfifo_produce <= 3'd0;
		soc_ethmac_crc32_checker_syncfifo_consume <= 3'd0;
		soc_ethmac_rx_converter_converter_source_first <= 1'd0;
		soc_ethmac_rx_converter_converter_source_last <= 1'd0;
		soc_ethmac_rx_converter_converter_demux <= 2'd0;
		soc_ethmac_rx_converter_converter_strobe_all <= 1'd0;
		soc_ethmac_rx_cdc_graycounter0_q <= 7'd0;
		soc_ethmac_rx_cdc_graycounter0_q_binary <= 7'd0;
		vns_clockdomainsrenamer1_state <= 1'd0;
		vns_clockdomainsrenamer3_state <= 2'd0;
		vns_clockdomainsrenamer5_state <= 2'd0;
	end
	vns_xilinxmultiregimpl5_regs0 <= soc_ethmac_rx_cdc_graycounter1_q;
	vns_xilinxmultiregimpl5_regs1 <= vns_xilinxmultiregimpl5_regs0;
end

always @(posedge eth_tx_clk) begin
	if (soc_ethmac_tx_gap_inserter_counter_reset) begin
		soc_ethmac_tx_gap_inserter_counter <= 1'd0;
	end else begin
		if (soc_ethmac_tx_gap_inserter_counter_ce) begin
			soc_ethmac_tx_gap_inserter_counter <= (soc_ethmac_tx_gap_inserter_counter + 1'd1);
		end
	end
	vns_clockdomainsrenamer0_state <= vns_clockdomainsrenamer0_next_state;
	if (soc_ethmac_preamble_inserter_clr_cnt) begin
		soc_ethmac_preamble_inserter_cnt <= 1'd0;
	end else begin
		if (soc_ethmac_preamble_inserter_inc_cnt) begin
			soc_ethmac_preamble_inserter_cnt <= (soc_ethmac_preamble_inserter_cnt + 1'd1);
		end
	end
	vns_clockdomainsrenamer2_state <= vns_clockdomainsrenamer2_next_state;
	if (soc_ethmac_crc32_inserter_is_ongoing0) begin
		soc_ethmac_crc32_inserter_cnt <= 2'd3;
	end else begin
		if ((soc_ethmac_crc32_inserter_is_ongoing1 & (~soc_ethmac_crc32_inserter_cnt_done))) begin
			soc_ethmac_crc32_inserter_cnt <= (soc_ethmac_crc32_inserter_cnt - soc_ethmac_crc32_inserter_source_ready);
		end
	end
	if (soc_ethmac_crc32_inserter_ce) begin
		soc_ethmac_crc32_inserter_reg <= soc_ethmac_crc32_inserter_next;
	end
	if (soc_ethmac_crc32_inserter_reset) begin
		soc_ethmac_crc32_inserter_reg <= 32'd4294967295;
	end
	vns_clockdomainsrenamer4_state <= vns_clockdomainsrenamer4_next_state;
	if (soc_ethmac_padding_inserter_counter_reset) begin
		soc_ethmac_padding_inserter_counter <= 1'd0;
	end else begin
		if (soc_ethmac_padding_inserter_counter_ce) begin
			soc_ethmac_padding_inserter_counter <= (soc_ethmac_padding_inserter_counter + 1'd1);
		end
	end
	vns_clockdomainsrenamer6_state <= vns_clockdomainsrenamer6_next_state;
	if ((soc_ethmac_tx_last_be_sink_valid & soc_ethmac_tx_last_be_sink_ready)) begin
		if (soc_ethmac_tx_last_be_sink_last) begin
			soc_ethmac_tx_last_be_ongoing <= 1'd1;
		end else begin
			if (soc_ethmac_tx_last_be_sink_payload_last_be) begin
				soc_ethmac_tx_last_be_ongoing <= 1'd0;
			end
		end
	end
	if ((soc_ethmac_tx_converter_converter_source_valid & soc_ethmac_tx_converter_converter_source_ready)) begin
		if (soc_ethmac_tx_converter_converter_last) begin
			soc_ethmac_tx_converter_converter_mux <= 1'd0;
		end else begin
			soc_ethmac_tx_converter_converter_mux <= (soc_ethmac_tx_converter_converter_mux + 1'd1);
		end
	end
	soc_ethmac_tx_cdc_graycounter1_q_binary <= soc_ethmac_tx_cdc_graycounter1_q_next_binary;
	soc_ethmac_tx_cdc_graycounter1_q <= soc_ethmac_tx_cdc_graycounter1_q_next;
	if (eth_tx_rst) begin
		soc_ethmac_crc32_inserter_reg <= 32'd4294967295;
		soc_ethmac_crc32_inserter_cnt <= 2'd3;
		soc_ethmac_padding_inserter_counter <= 16'd1;
		soc_ethmac_tx_last_be_ongoing <= 1'd1;
		soc_ethmac_tx_converter_converter_mux <= 2'd0;
		soc_ethmac_tx_cdc_graycounter1_q <= 7'd0;
		soc_ethmac_tx_cdc_graycounter1_q_binary <= 7'd0;
		vns_clockdomainsrenamer0_state <= 1'd0;
		vns_clockdomainsrenamer2_state <= 2'd0;
		vns_clockdomainsrenamer4_state <= 2'd0;
		vns_clockdomainsrenamer6_state <= 1'd0;
	end
	vns_xilinxmultiregimpl2_regs0 <= soc_ethmac_tx_cdc_graycounter0_q;
	vns_xilinxmultiregimpl2_regs1 <= vns_xilinxmultiregimpl2_regs0;
end

always @(posedge fmeter_clk) begin
	soc_hdmi_in0_freq_q_binary <= soc_hdmi_in0_freq_q_next_binary;
	soc_hdmi_in0_freq_q <= soc_hdmi_in0_freq_q_next;
end

always @(posedge hdmi_in0_pix_clk) begin
	soc_charsync0_raw_data1 <= soc_charsync0_raw_data;
	soc_charsync0_found_control <= 1'd0;
	if (((((soc_charsync0_raw[9:0] == 10'd852) | (soc_charsync0_raw[9:0] == 8'd171)) | (soc_charsync0_raw[9:0] == 9'd340)) | (soc_charsync0_raw[9:0] == 10'd683))) begin
		soc_charsync0_found_control <= 1'd1;
		soc_charsync0_control_position <= 1'd0;
	end
	if (((((soc_charsync0_raw[10:1] == 10'd852) | (soc_charsync0_raw[10:1] == 8'd171)) | (soc_charsync0_raw[10:1] == 9'd340)) | (soc_charsync0_raw[10:1] == 10'd683))) begin
		soc_charsync0_found_control <= 1'd1;
		soc_charsync0_control_position <= 1'd1;
	end
	if (((((soc_charsync0_raw[11:2] == 10'd852) | (soc_charsync0_raw[11:2] == 8'd171)) | (soc_charsync0_raw[11:2] == 9'd340)) | (soc_charsync0_raw[11:2] == 10'd683))) begin
		soc_charsync0_found_control <= 1'd1;
		soc_charsync0_control_position <= 2'd2;
	end
	if (((((soc_charsync0_raw[12:3] == 10'd852) | (soc_charsync0_raw[12:3] == 8'd171)) | (soc_charsync0_raw[12:3] == 9'd340)) | (soc_charsync0_raw[12:3] == 10'd683))) begin
		soc_charsync0_found_control <= 1'd1;
		soc_charsync0_control_position <= 2'd3;
	end
	if (((((soc_charsync0_raw[13:4] == 10'd852) | (soc_charsync0_raw[13:4] == 8'd171)) | (soc_charsync0_raw[13:4] == 9'd340)) | (soc_charsync0_raw[13:4] == 10'd683))) begin
		soc_charsync0_found_control <= 1'd1;
		soc_charsync0_control_position <= 3'd4;
	end
	if (((((soc_charsync0_raw[14:5] == 10'd852) | (soc_charsync0_raw[14:5] == 8'd171)) | (soc_charsync0_raw[14:5] == 9'd340)) | (soc_charsync0_raw[14:5] == 10'd683))) begin
		soc_charsync0_found_control <= 1'd1;
		soc_charsync0_control_position <= 3'd5;
	end
	if (((((soc_charsync0_raw[15:6] == 10'd852) | (soc_charsync0_raw[15:6] == 8'd171)) | (soc_charsync0_raw[15:6] == 9'd340)) | (soc_charsync0_raw[15:6] == 10'd683))) begin
		soc_charsync0_found_control <= 1'd1;
		soc_charsync0_control_position <= 3'd6;
	end
	if (((((soc_charsync0_raw[16:7] == 10'd852) | (soc_charsync0_raw[16:7] == 8'd171)) | (soc_charsync0_raw[16:7] == 9'd340)) | (soc_charsync0_raw[16:7] == 10'd683))) begin
		soc_charsync0_found_control <= 1'd1;
		soc_charsync0_control_position <= 3'd7;
	end
	if (((((soc_charsync0_raw[17:8] == 10'd852) | (soc_charsync0_raw[17:8] == 8'd171)) | (soc_charsync0_raw[17:8] == 9'd340)) | (soc_charsync0_raw[17:8] == 10'd683))) begin
		soc_charsync0_found_control <= 1'd1;
		soc_charsync0_control_position <= 4'd8;
	end
	if (((((soc_charsync0_raw[18:9] == 10'd852) | (soc_charsync0_raw[18:9] == 8'd171)) | (soc_charsync0_raw[18:9] == 9'd340)) | (soc_charsync0_raw[18:9] == 10'd683))) begin
		soc_charsync0_found_control <= 1'd1;
		soc_charsync0_control_position <= 4'd9;
	end
	if ((soc_charsync0_found_control & (soc_charsync0_control_position == soc_charsync0_previous_control_position))) begin
		if ((soc_charsync0_control_counter == 3'd7)) begin
			soc_charsync0_control_counter <= 1'd0;
			soc_charsync0_synced <= 1'd1;
			soc_charsync0_word_sel <= soc_charsync0_control_position;
		end else begin
			soc_charsync0_control_counter <= (soc_charsync0_control_counter + 1'd1);
		end
	end else begin
		soc_charsync0_control_counter <= 1'd0;
	end
	soc_charsync0_previous_control_position <= soc_charsync0_control_position;
	soc_charsync0_data <= (soc_charsync0_raw >>> soc_charsync0_word_sel);
	soc_wer0_data_r <= soc_wer0_data[8:0];
	soc_wer0_transition_count <= (((((((soc_wer0_transitions[0] + soc_wer0_transitions[1]) + soc_wer0_transitions[2]) + soc_wer0_transitions[3]) + soc_wer0_transitions[4]) + soc_wer0_transitions[5]) + soc_wer0_transitions[6]) + soc_wer0_transitions[7]);
	soc_wer0_is_control <= ((((soc_wer0_data_r == 10'd852) | (soc_wer0_data_r == 8'd171)) | (soc_wer0_data_r == 9'd340)) | (soc_wer0_data_r == 10'd683));
	soc_wer0_is_error <= ((soc_wer0_transition_count > 3'd4) & (~soc_wer0_is_control));
	{soc_wer0_period_done, soc_wer0_period_counter} <= (soc_wer0_period_counter + 1'd1);
	soc_wer0_wer_counter_r_updated <= soc_wer0_period_done;
	if (soc_wer0_period_done) begin
		soc_wer0_wer_counter_r <= soc_wer0_wer_counter;
		soc_wer0_wer_counter <= 1'd0;
	end else begin
		if (soc_wer0_is_error) begin
			soc_wer0_wer_counter <= (soc_wer0_wer_counter + 1'd1);
		end
	end
	if (soc_wer0_i) begin
		soc_wer0_toggle_i <= (~soc_wer0_toggle_i);
	end
	soc_decoding0_output_de <= 1'd1;
	if ((soc_decoding0_input == 10'd852)) begin
		soc_decoding0_output_de <= 1'd0;
		soc_decoding0_output_c <= 1'd0;
	end
	if ((soc_decoding0_input == 8'd171)) begin
		soc_decoding0_output_de <= 1'd0;
		soc_decoding0_output_c <= 1'd1;
	end
	if ((soc_decoding0_input == 9'd340)) begin
		soc_decoding0_output_de <= 1'd0;
		soc_decoding0_output_c <= 2'd2;
	end
	if ((soc_decoding0_input == 10'd683)) begin
		soc_decoding0_output_de <= 1'd0;
		soc_decoding0_output_c <= 2'd3;
	end
	soc_decoding0_output_d[0] <= (soc_decoding0_input[0] ^ soc_decoding0_input[9]);
	soc_decoding0_output_d[1] <= ((soc_decoding0_input[1] ^ soc_decoding0_input[0]) ^ (~soc_decoding0_input[8]));
	soc_decoding0_output_d[2] <= ((soc_decoding0_input[2] ^ soc_decoding0_input[1]) ^ (~soc_decoding0_input[8]));
	soc_decoding0_output_d[3] <= ((soc_decoding0_input[3] ^ soc_decoding0_input[2]) ^ (~soc_decoding0_input[8]));
	soc_decoding0_output_d[4] <= ((soc_decoding0_input[4] ^ soc_decoding0_input[3]) ^ (~soc_decoding0_input[8]));
	soc_decoding0_output_d[5] <= ((soc_decoding0_input[5] ^ soc_decoding0_input[4]) ^ (~soc_decoding0_input[8]));
	soc_decoding0_output_d[6] <= ((soc_decoding0_input[6] ^ soc_decoding0_input[5]) ^ (~soc_decoding0_input[8]));
	soc_decoding0_output_d[7] <= ((soc_decoding0_input[7] ^ soc_decoding0_input[6]) ^ (~soc_decoding0_input[8]));
	soc_decoding0_valid_o <= soc_decoding0_valid_i;
	soc_charsync1_raw_data1 <= soc_charsync1_raw_data;
	soc_charsync1_found_control <= 1'd0;
	if (((((soc_charsync1_raw[9:0] == 10'd852) | (soc_charsync1_raw[9:0] == 8'd171)) | (soc_charsync1_raw[9:0] == 9'd340)) | (soc_charsync1_raw[9:0] == 10'd683))) begin
		soc_charsync1_found_control <= 1'd1;
		soc_charsync1_control_position <= 1'd0;
	end
	if (((((soc_charsync1_raw[10:1] == 10'd852) | (soc_charsync1_raw[10:1] == 8'd171)) | (soc_charsync1_raw[10:1] == 9'd340)) | (soc_charsync1_raw[10:1] == 10'd683))) begin
		soc_charsync1_found_control <= 1'd1;
		soc_charsync1_control_position <= 1'd1;
	end
	if (((((soc_charsync1_raw[11:2] == 10'd852) | (soc_charsync1_raw[11:2] == 8'd171)) | (soc_charsync1_raw[11:2] == 9'd340)) | (soc_charsync1_raw[11:2] == 10'd683))) begin
		soc_charsync1_found_control <= 1'd1;
		soc_charsync1_control_position <= 2'd2;
	end
	if (((((soc_charsync1_raw[12:3] == 10'd852) | (soc_charsync1_raw[12:3] == 8'd171)) | (soc_charsync1_raw[12:3] == 9'd340)) | (soc_charsync1_raw[12:3] == 10'd683))) begin
		soc_charsync1_found_control <= 1'd1;
		soc_charsync1_control_position <= 2'd3;
	end
	if (((((soc_charsync1_raw[13:4] == 10'd852) | (soc_charsync1_raw[13:4] == 8'd171)) | (soc_charsync1_raw[13:4] == 9'd340)) | (soc_charsync1_raw[13:4] == 10'd683))) begin
		soc_charsync1_found_control <= 1'd1;
		soc_charsync1_control_position <= 3'd4;
	end
	if (((((soc_charsync1_raw[14:5] == 10'd852) | (soc_charsync1_raw[14:5] == 8'd171)) | (soc_charsync1_raw[14:5] == 9'd340)) | (soc_charsync1_raw[14:5] == 10'd683))) begin
		soc_charsync1_found_control <= 1'd1;
		soc_charsync1_control_position <= 3'd5;
	end
	if (((((soc_charsync1_raw[15:6] == 10'd852) | (soc_charsync1_raw[15:6] == 8'd171)) | (soc_charsync1_raw[15:6] == 9'd340)) | (soc_charsync1_raw[15:6] == 10'd683))) begin
		soc_charsync1_found_control <= 1'd1;
		soc_charsync1_control_position <= 3'd6;
	end
	if (((((soc_charsync1_raw[16:7] == 10'd852) | (soc_charsync1_raw[16:7] == 8'd171)) | (soc_charsync1_raw[16:7] == 9'd340)) | (soc_charsync1_raw[16:7] == 10'd683))) begin
		soc_charsync1_found_control <= 1'd1;
		soc_charsync1_control_position <= 3'd7;
	end
	if (((((soc_charsync1_raw[17:8] == 10'd852) | (soc_charsync1_raw[17:8] == 8'd171)) | (soc_charsync1_raw[17:8] == 9'd340)) | (soc_charsync1_raw[17:8] == 10'd683))) begin
		soc_charsync1_found_control <= 1'd1;
		soc_charsync1_control_position <= 4'd8;
	end
	if (((((soc_charsync1_raw[18:9] == 10'd852) | (soc_charsync1_raw[18:9] == 8'd171)) | (soc_charsync1_raw[18:9] == 9'd340)) | (soc_charsync1_raw[18:9] == 10'd683))) begin
		soc_charsync1_found_control <= 1'd1;
		soc_charsync1_control_position <= 4'd9;
	end
	if ((soc_charsync1_found_control & (soc_charsync1_control_position == soc_charsync1_previous_control_position))) begin
		if ((soc_charsync1_control_counter == 3'd7)) begin
			soc_charsync1_control_counter <= 1'd0;
			soc_charsync1_synced <= 1'd1;
			soc_charsync1_word_sel <= soc_charsync1_control_position;
		end else begin
			soc_charsync1_control_counter <= (soc_charsync1_control_counter + 1'd1);
		end
	end else begin
		soc_charsync1_control_counter <= 1'd0;
	end
	soc_charsync1_previous_control_position <= soc_charsync1_control_position;
	soc_charsync1_data <= (soc_charsync1_raw >>> soc_charsync1_word_sel);
	soc_wer1_data_r <= soc_wer1_data[8:0];
	soc_wer1_transition_count <= (((((((soc_wer1_transitions[0] + soc_wer1_transitions[1]) + soc_wer1_transitions[2]) + soc_wer1_transitions[3]) + soc_wer1_transitions[4]) + soc_wer1_transitions[5]) + soc_wer1_transitions[6]) + soc_wer1_transitions[7]);
	soc_wer1_is_control <= ((((soc_wer1_data_r == 10'd852) | (soc_wer1_data_r == 8'd171)) | (soc_wer1_data_r == 9'd340)) | (soc_wer1_data_r == 10'd683));
	soc_wer1_is_error <= ((soc_wer1_transition_count > 3'd4) & (~soc_wer1_is_control));
	{soc_wer1_period_done, soc_wer1_period_counter} <= (soc_wer1_period_counter + 1'd1);
	soc_wer1_wer_counter_r_updated <= soc_wer1_period_done;
	if (soc_wer1_period_done) begin
		soc_wer1_wer_counter_r <= soc_wer1_wer_counter;
		soc_wer1_wer_counter <= 1'd0;
	end else begin
		if (soc_wer1_is_error) begin
			soc_wer1_wer_counter <= (soc_wer1_wer_counter + 1'd1);
		end
	end
	if (soc_wer1_i) begin
		soc_wer1_toggle_i <= (~soc_wer1_toggle_i);
	end
	soc_decoding1_output_de <= 1'd1;
	if ((soc_decoding1_input == 10'd852)) begin
		soc_decoding1_output_de <= 1'd0;
		soc_decoding1_output_c <= 1'd0;
	end
	if ((soc_decoding1_input == 8'd171)) begin
		soc_decoding1_output_de <= 1'd0;
		soc_decoding1_output_c <= 1'd1;
	end
	if ((soc_decoding1_input == 9'd340)) begin
		soc_decoding1_output_de <= 1'd0;
		soc_decoding1_output_c <= 2'd2;
	end
	if ((soc_decoding1_input == 10'd683)) begin
		soc_decoding1_output_de <= 1'd0;
		soc_decoding1_output_c <= 2'd3;
	end
	soc_decoding1_output_d[0] <= (soc_decoding1_input[0] ^ soc_decoding1_input[9]);
	soc_decoding1_output_d[1] <= ((soc_decoding1_input[1] ^ soc_decoding1_input[0]) ^ (~soc_decoding1_input[8]));
	soc_decoding1_output_d[2] <= ((soc_decoding1_input[2] ^ soc_decoding1_input[1]) ^ (~soc_decoding1_input[8]));
	soc_decoding1_output_d[3] <= ((soc_decoding1_input[3] ^ soc_decoding1_input[2]) ^ (~soc_decoding1_input[8]));
	soc_decoding1_output_d[4] <= ((soc_decoding1_input[4] ^ soc_decoding1_input[3]) ^ (~soc_decoding1_input[8]));
	soc_decoding1_output_d[5] <= ((soc_decoding1_input[5] ^ soc_decoding1_input[4]) ^ (~soc_decoding1_input[8]));
	soc_decoding1_output_d[6] <= ((soc_decoding1_input[6] ^ soc_decoding1_input[5]) ^ (~soc_decoding1_input[8]));
	soc_decoding1_output_d[7] <= ((soc_decoding1_input[7] ^ soc_decoding1_input[6]) ^ (~soc_decoding1_input[8]));
	soc_decoding1_valid_o <= soc_decoding1_valid_i;
	soc_charsync2_raw_data1 <= soc_charsync2_raw_data;
	soc_charsync2_found_control <= 1'd0;
	if (((((soc_charsync2_raw[9:0] == 10'd852) | (soc_charsync2_raw[9:0] == 8'd171)) | (soc_charsync2_raw[9:0] == 9'd340)) | (soc_charsync2_raw[9:0] == 10'd683))) begin
		soc_charsync2_found_control <= 1'd1;
		soc_charsync2_control_position <= 1'd0;
	end
	if (((((soc_charsync2_raw[10:1] == 10'd852) | (soc_charsync2_raw[10:1] == 8'd171)) | (soc_charsync2_raw[10:1] == 9'd340)) | (soc_charsync2_raw[10:1] == 10'd683))) begin
		soc_charsync2_found_control <= 1'd1;
		soc_charsync2_control_position <= 1'd1;
	end
	if (((((soc_charsync2_raw[11:2] == 10'd852) | (soc_charsync2_raw[11:2] == 8'd171)) | (soc_charsync2_raw[11:2] == 9'd340)) | (soc_charsync2_raw[11:2] == 10'd683))) begin
		soc_charsync2_found_control <= 1'd1;
		soc_charsync2_control_position <= 2'd2;
	end
	if (((((soc_charsync2_raw[12:3] == 10'd852) | (soc_charsync2_raw[12:3] == 8'd171)) | (soc_charsync2_raw[12:3] == 9'd340)) | (soc_charsync2_raw[12:3] == 10'd683))) begin
		soc_charsync2_found_control <= 1'd1;
		soc_charsync2_control_position <= 2'd3;
	end
	if (((((soc_charsync2_raw[13:4] == 10'd852) | (soc_charsync2_raw[13:4] == 8'd171)) | (soc_charsync2_raw[13:4] == 9'd340)) | (soc_charsync2_raw[13:4] == 10'd683))) begin
		soc_charsync2_found_control <= 1'd1;
		soc_charsync2_control_position <= 3'd4;
	end
	if (((((soc_charsync2_raw[14:5] == 10'd852) | (soc_charsync2_raw[14:5] == 8'd171)) | (soc_charsync2_raw[14:5] == 9'd340)) | (soc_charsync2_raw[14:5] == 10'd683))) begin
		soc_charsync2_found_control <= 1'd1;
		soc_charsync2_control_position <= 3'd5;
	end
	if (((((soc_charsync2_raw[15:6] == 10'd852) | (soc_charsync2_raw[15:6] == 8'd171)) | (soc_charsync2_raw[15:6] == 9'd340)) | (soc_charsync2_raw[15:6] == 10'd683))) begin
		soc_charsync2_found_control <= 1'd1;
		soc_charsync2_control_position <= 3'd6;
	end
	if (((((soc_charsync2_raw[16:7] == 10'd852) | (soc_charsync2_raw[16:7] == 8'd171)) | (soc_charsync2_raw[16:7] == 9'd340)) | (soc_charsync2_raw[16:7] == 10'd683))) begin
		soc_charsync2_found_control <= 1'd1;
		soc_charsync2_control_position <= 3'd7;
	end
	if (((((soc_charsync2_raw[17:8] == 10'd852) | (soc_charsync2_raw[17:8] == 8'd171)) | (soc_charsync2_raw[17:8] == 9'd340)) | (soc_charsync2_raw[17:8] == 10'd683))) begin
		soc_charsync2_found_control <= 1'd1;
		soc_charsync2_control_position <= 4'd8;
	end
	if (((((soc_charsync2_raw[18:9] == 10'd852) | (soc_charsync2_raw[18:9] == 8'd171)) | (soc_charsync2_raw[18:9] == 9'd340)) | (soc_charsync2_raw[18:9] == 10'd683))) begin
		soc_charsync2_found_control <= 1'd1;
		soc_charsync2_control_position <= 4'd9;
	end
	if ((soc_charsync2_found_control & (soc_charsync2_control_position == soc_charsync2_previous_control_position))) begin
		if ((soc_charsync2_control_counter == 3'd7)) begin
			soc_charsync2_control_counter <= 1'd0;
			soc_charsync2_synced <= 1'd1;
			soc_charsync2_word_sel <= soc_charsync2_control_position;
		end else begin
			soc_charsync2_control_counter <= (soc_charsync2_control_counter + 1'd1);
		end
	end else begin
		soc_charsync2_control_counter <= 1'd0;
	end
	soc_charsync2_previous_control_position <= soc_charsync2_control_position;
	soc_charsync2_data <= (soc_charsync2_raw >>> soc_charsync2_word_sel);
	soc_wer2_data_r <= soc_wer2_data[8:0];
	soc_wer2_transition_count <= (((((((soc_wer2_transitions[0] + soc_wer2_transitions[1]) + soc_wer2_transitions[2]) + soc_wer2_transitions[3]) + soc_wer2_transitions[4]) + soc_wer2_transitions[5]) + soc_wer2_transitions[6]) + soc_wer2_transitions[7]);
	soc_wer2_is_control <= ((((soc_wer2_data_r == 10'd852) | (soc_wer2_data_r == 8'd171)) | (soc_wer2_data_r == 9'd340)) | (soc_wer2_data_r == 10'd683));
	soc_wer2_is_error <= ((soc_wer2_transition_count > 3'd4) & (~soc_wer2_is_control));
	{soc_wer2_period_done, soc_wer2_period_counter} <= (soc_wer2_period_counter + 1'd1);
	soc_wer2_wer_counter_r_updated <= soc_wer2_period_done;
	if (soc_wer2_period_done) begin
		soc_wer2_wer_counter_r <= soc_wer2_wer_counter;
		soc_wer2_wer_counter <= 1'd0;
	end else begin
		if (soc_wer2_is_error) begin
			soc_wer2_wer_counter <= (soc_wer2_wer_counter + 1'd1);
		end
	end
	if (soc_wer2_i) begin
		soc_wer2_toggle_i <= (~soc_wer2_toggle_i);
	end
	soc_decoding2_output_de <= 1'd1;
	if ((soc_decoding2_input == 10'd852)) begin
		soc_decoding2_output_de <= 1'd0;
		soc_decoding2_output_c <= 1'd0;
	end
	if ((soc_decoding2_input == 8'd171)) begin
		soc_decoding2_output_de <= 1'd0;
		soc_decoding2_output_c <= 1'd1;
	end
	if ((soc_decoding2_input == 9'd340)) begin
		soc_decoding2_output_de <= 1'd0;
		soc_decoding2_output_c <= 2'd2;
	end
	if ((soc_decoding2_input == 10'd683)) begin
		soc_decoding2_output_de <= 1'd0;
		soc_decoding2_output_c <= 2'd3;
	end
	soc_decoding2_output_d[0] <= (soc_decoding2_input[0] ^ soc_decoding2_input[9]);
	soc_decoding2_output_d[1] <= ((soc_decoding2_input[1] ^ soc_decoding2_input[0]) ^ (~soc_decoding2_input[8]));
	soc_decoding2_output_d[2] <= ((soc_decoding2_input[2] ^ soc_decoding2_input[1]) ^ (~soc_decoding2_input[8]));
	soc_decoding2_output_d[3] <= ((soc_decoding2_input[3] ^ soc_decoding2_input[2]) ^ (~soc_decoding2_input[8]));
	soc_decoding2_output_d[4] <= ((soc_decoding2_input[4] ^ soc_decoding2_input[3]) ^ (~soc_decoding2_input[8]));
	soc_decoding2_output_d[5] <= ((soc_decoding2_input[5] ^ soc_decoding2_input[4]) ^ (~soc_decoding2_input[8]));
	soc_decoding2_output_d[6] <= ((soc_decoding2_input[6] ^ soc_decoding2_input[5]) ^ (~soc_decoding2_input[8]));
	soc_decoding2_output_d[7] <= ((soc_decoding2_input[7] ^ soc_decoding2_input[6]) ^ (~soc_decoding2_input[8]));
	soc_decoding2_valid_o <= soc_decoding2_valid_i;
	if ((~soc_chansync_valid_i)) begin
		soc_chansync_chan_synced <= 1'd0;
	end else begin
		if (soc_chansync_some_control) begin
			if (soc_chansync_all_control) begin
				soc_chansync_chan_synced <= 1'd1;
			end else begin
				soc_chansync_chan_synced <= 1'd0;
			end
		end
	end
	soc_chansync_syncbuffer0_produce <= (soc_chansync_syncbuffer0_produce + 1'd1);
	if (soc_chansync_syncbuffer0_re) begin
		soc_chansync_syncbuffer0_consume <= (soc_chansync_syncbuffer0_consume + 1'd1);
	end
	soc_chansync_syncbuffer1_produce <= (soc_chansync_syncbuffer1_produce + 1'd1);
	if (soc_chansync_syncbuffer1_re) begin
		soc_chansync_syncbuffer1_consume <= (soc_chansync_syncbuffer1_consume + 1'd1);
	end
	soc_chansync_syncbuffer2_produce <= (soc_chansync_syncbuffer2_produce + 1'd1);
	if (soc_chansync_syncbuffer2_re) begin
		soc_chansync_syncbuffer2_consume <= (soc_chansync_syncbuffer2_consume + 1'd1);
	end
	soc_syncpol_valid_o <= soc_syncpol_valid_i;
	soc_syncpol_r <= soc_syncpol_data_in2_d;
	soc_syncpol_g <= soc_syncpol_data_in1_d;
	soc_syncpol_b <= soc_syncpol_data_in0_d;
	soc_syncpol_de_r <= soc_syncpol_data_in0_de;
	if ((soc_syncpol_de_r & (~soc_syncpol_data_in0_de))) begin
		soc_syncpol_c_polarity <= soc_syncpol_data_in0_c;
		soc_syncpol_c_out <= 1'd0;
	end else begin
		soc_syncpol_c_out <= (soc_syncpol_data_in0_c ^ soc_syncpol_c_polarity);
	end
	soc_resdetection_de_r <= soc_resdetection_de;
	if ((soc_resdetection_valid_i & soc_resdetection_de)) begin
		soc_resdetection_hcounter <= (soc_resdetection_hcounter + 1'd1);
	end else begin
		soc_resdetection_hcounter <= 1'd0;
	end
	if (soc_resdetection_valid_i) begin
		if (soc_resdetection_pn_de) begin
			soc_resdetection_hcounter_st <= soc_resdetection_hcounter;
		end
	end else begin
		soc_resdetection_hcounter_st <= 1'd0;
	end
	soc_resdetection_vsync_r <= soc_resdetection_vsync;
	if ((soc_resdetection_valid_i & soc_resdetection_p_vsync)) begin
		soc_resdetection_vcounter <= 1'd0;
	end else begin
		if (soc_resdetection_pn_de) begin
			soc_resdetection_vcounter <= (soc_resdetection_vcounter + 1'd1);
		end
	end
	if (soc_resdetection_valid_i) begin
		if (soc_resdetection_p_vsync) begin
			soc_resdetection_vcounter_st <= soc_resdetection_vcounter;
		end
	end else begin
		soc_resdetection_vcounter_st <= 1'd0;
	end
	soc_frame_de_r <= soc_frame_de;
	soc_frame_next_de0 <= soc_frame_de;
	soc_frame_next_vsync0 <= soc_frame_vsync;
	soc_frame_next_de1 <= soc_frame_next_de0;
	soc_frame_next_vsync1 <= soc_frame_next_vsync0;
	soc_frame_next_de2 <= soc_frame_next_de1;
	soc_frame_next_vsync2 <= soc_frame_next_vsync1;
	soc_frame_next_de3 <= soc_frame_next_de2;
	soc_frame_next_vsync3 <= soc_frame_next_vsync2;
	soc_frame_next_de4 <= soc_frame_next_de3;
	soc_frame_next_vsync4 <= soc_frame_next_vsync3;
	soc_frame_next_de5 <= soc_frame_next_de4;
	soc_frame_next_vsync5 <= soc_frame_next_vsync4;
	soc_frame_next_de6 <= soc_frame_next_de5;
	soc_frame_next_vsync6 <= soc_frame_next_vsync5;
	soc_frame_next_de7 <= soc_frame_next_de6;
	soc_frame_next_vsync7 <= soc_frame_next_vsync6;
	soc_frame_next_de8 <= soc_frame_next_de7;
	soc_frame_next_vsync8 <= soc_frame_next_vsync7;
	soc_frame_next_de9 <= soc_frame_next_de8;
	soc_frame_next_vsync9 <= soc_frame_next_vsync8;
	soc_frame_next_de10 <= soc_frame_next_de9;
	soc_frame_next_vsync10 <= soc_frame_next_vsync9;
	soc_frame_vsync_r <= soc_frame_next_vsync10;
	soc_frame_cur_word_valid <= 1'd0;
	if (soc_frame_new_frame) begin
		soc_frame_cur_word_valid <= (soc_frame_pack_counter == 3'd7);
		soc_frame_pack_counter <= 1'd0;
	end else begin
		if ((soc_frame_chroma_downsampler_source_valid & soc_frame_next_de10)) begin
			if ((soc_frame_pack_counter == 3'd7)) begin
				soc_frame_cur_word[15:0] <= soc_frame_encoded_pixel;
			end
			if ((soc_frame_pack_counter == 3'd6)) begin
				soc_frame_cur_word[31:16] <= soc_frame_encoded_pixel;
			end
			if ((soc_frame_pack_counter == 3'd5)) begin
				soc_frame_cur_word[47:32] <= soc_frame_encoded_pixel;
			end
			if ((soc_frame_pack_counter == 3'd4)) begin
				soc_frame_cur_word[63:48] <= soc_frame_encoded_pixel;
			end
			if ((soc_frame_pack_counter == 2'd3)) begin
				soc_frame_cur_word[79:64] <= soc_frame_encoded_pixel;
			end
			if ((soc_frame_pack_counter == 2'd2)) begin
				soc_frame_cur_word[95:80] <= soc_frame_encoded_pixel;
			end
			if ((soc_frame_pack_counter == 1'd1)) begin
				soc_frame_cur_word[111:96] <= soc_frame_encoded_pixel;
			end
			if ((soc_frame_pack_counter == 1'd0)) begin
				soc_frame_cur_word[127:112] <= soc_frame_encoded_pixel;
			end
			soc_frame_cur_word_valid <= (soc_frame_pack_counter == 3'd7);
			soc_frame_pack_counter <= (soc_frame_pack_counter + 1'd1);
		end
	end
	if (soc_frame_new_frame) begin
		soc_frame_fifo_sink_payload_sof <= 1'd1;
	end else begin
		if (soc_frame_cur_word_valid) begin
			soc_frame_fifo_sink_payload_sof <= 1'd0;
		end
	end
	if ((soc_frame_fifo_sink_valid & (~soc_frame_fifo_sink_ready))) begin
		soc_frame_pix_overflow <= 1'd1;
	end else begin
		if (soc_frame_pix_overflow_reset) begin
			soc_frame_pix_overflow <= 1'd0;
		end
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_valid_n0 <= soc_frame_rgb2ycbcr_sink_valid;
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_valid_n1 <= soc_frame_rgb2ycbcr_valid_n0;
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_valid_n2 <= soc_frame_rgb2ycbcr_valid_n1;
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_valid_n3 <= soc_frame_rgb2ycbcr_valid_n2;
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_valid_n4 <= soc_frame_rgb2ycbcr_valid_n3;
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_valid_n5 <= soc_frame_rgb2ycbcr_valid_n4;
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_valid_n6 <= soc_frame_rgb2ycbcr_valid_n5;
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_valid_n7 <= soc_frame_rgb2ycbcr_valid_n6;
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_first_n0 <= (soc_frame_rgb2ycbcr_sink_valid & soc_frame_rgb2ycbcr_sink_first);
		soc_frame_rgb2ycbcr_last_n0 <= (soc_frame_rgb2ycbcr_sink_valid & soc_frame_rgb2ycbcr_sink_last);
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_first_n1 <= soc_frame_rgb2ycbcr_first_n0;
		soc_frame_rgb2ycbcr_last_n1 <= soc_frame_rgb2ycbcr_last_n0;
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_first_n2 <= soc_frame_rgb2ycbcr_first_n1;
		soc_frame_rgb2ycbcr_last_n2 <= soc_frame_rgb2ycbcr_last_n1;
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_first_n3 <= soc_frame_rgb2ycbcr_first_n2;
		soc_frame_rgb2ycbcr_last_n3 <= soc_frame_rgb2ycbcr_last_n2;
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_first_n4 <= soc_frame_rgb2ycbcr_first_n3;
		soc_frame_rgb2ycbcr_last_n4 <= soc_frame_rgb2ycbcr_last_n3;
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_first_n5 <= soc_frame_rgb2ycbcr_first_n4;
		soc_frame_rgb2ycbcr_last_n5 <= soc_frame_rgb2ycbcr_last_n4;
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_first_n6 <= soc_frame_rgb2ycbcr_first_n5;
		soc_frame_rgb2ycbcr_last_n6 <= soc_frame_rgb2ycbcr_last_n5;
	end
	if (soc_frame_rgb2ycbcr_pipe_ce) begin
		soc_frame_rgb2ycbcr_first_n7 <= soc_frame_rgb2ycbcr_first_n6;
		soc_frame_rgb2ycbcr_last_n7 <= soc_frame_rgb2ycbcr_last_n6;
	end
	if (soc_frame_rgb2ycbcr_ce) begin
		soc_frame_rgb2ycbcr_record0_rgb_n_r <= soc_frame_rgb2ycbcr_sink_r;
		soc_frame_rgb2ycbcr_record0_rgb_n_g <= soc_frame_rgb2ycbcr_sink_g;
		soc_frame_rgb2ycbcr_record0_rgb_n_b <= soc_frame_rgb2ycbcr_sink_b;
		soc_frame_rgb2ycbcr_record1_rgb_n_r <= soc_frame_rgb2ycbcr_record0_rgb_n_r;
		soc_frame_rgb2ycbcr_record1_rgb_n_g <= soc_frame_rgb2ycbcr_record0_rgb_n_g;
		soc_frame_rgb2ycbcr_record1_rgb_n_b <= soc_frame_rgb2ycbcr_record0_rgb_n_b;
		soc_frame_rgb2ycbcr_record2_rgb_n_r <= soc_frame_rgb2ycbcr_record1_rgb_n_r;
		soc_frame_rgb2ycbcr_record2_rgb_n_g <= soc_frame_rgb2ycbcr_record1_rgb_n_g;
		soc_frame_rgb2ycbcr_record2_rgb_n_b <= soc_frame_rgb2ycbcr_record1_rgb_n_b;
		soc_frame_rgb2ycbcr_record3_rgb_n_r <= soc_frame_rgb2ycbcr_record2_rgb_n_r;
		soc_frame_rgb2ycbcr_record3_rgb_n_g <= soc_frame_rgb2ycbcr_record2_rgb_n_g;
		soc_frame_rgb2ycbcr_record3_rgb_n_b <= soc_frame_rgb2ycbcr_record2_rgb_n_b;
		soc_frame_rgb2ycbcr_record4_rgb_n_r <= soc_frame_rgb2ycbcr_record3_rgb_n_r;
		soc_frame_rgb2ycbcr_record4_rgb_n_g <= soc_frame_rgb2ycbcr_record3_rgb_n_g;
		soc_frame_rgb2ycbcr_record4_rgb_n_b <= soc_frame_rgb2ycbcr_record3_rgb_n_b;
		soc_frame_rgb2ycbcr_record5_rgb_n_r <= soc_frame_rgb2ycbcr_record4_rgb_n_r;
		soc_frame_rgb2ycbcr_record5_rgb_n_g <= soc_frame_rgb2ycbcr_record4_rgb_n_g;
		soc_frame_rgb2ycbcr_record5_rgb_n_b <= soc_frame_rgb2ycbcr_record4_rgb_n_b;
		soc_frame_rgb2ycbcr_record6_rgb_n_r <= soc_frame_rgb2ycbcr_record5_rgb_n_r;
		soc_frame_rgb2ycbcr_record6_rgb_n_g <= soc_frame_rgb2ycbcr_record5_rgb_n_g;
		soc_frame_rgb2ycbcr_record6_rgb_n_b <= soc_frame_rgb2ycbcr_record5_rgb_n_b;
		soc_frame_rgb2ycbcr_record7_rgb_n_r <= soc_frame_rgb2ycbcr_record6_rgb_n_r;
		soc_frame_rgb2ycbcr_record7_rgb_n_g <= soc_frame_rgb2ycbcr_record6_rgb_n_g;
		soc_frame_rgb2ycbcr_record7_rgb_n_b <= soc_frame_rgb2ycbcr_record6_rgb_n_b;
		soc_frame_rgb2ycbcr_r_minus_g <= (soc_frame_rgb2ycbcr_sink_r - soc_frame_rgb2ycbcr_sink_g);
		soc_frame_rgb2ycbcr_b_minus_g <= (soc_frame_rgb2ycbcr_sink_b - soc_frame_rgb2ycbcr_sink_g);
		soc_frame_rgb2ycbcr_ca_mult_rg <= (soc_frame_rgb2ycbcr_r_minus_g * $signed({1'd0, 6'd46}));
		soc_frame_rgb2ycbcr_cb_mult_bg <= (soc_frame_rgb2ycbcr_b_minus_g * $signed({1'd0, 4'd15}));
		soc_frame_rgb2ycbcr_carg_plus_cbbg <= (soc_frame_rgb2ycbcr_ca_mult_rg + soc_frame_rgb2ycbcr_cb_mult_bg);
		soc_frame_rgb2ycbcr_yraw <= (soc_frame_rgb2ycbcr_carg_plus_cbbg[24:8] + $signed({1'd0, soc_frame_rgb2ycbcr_record2_rgb_n_g}));
		soc_frame_rgb2ycbcr_b_minus_yraw <= ($signed({1'd0, soc_frame_rgb2ycbcr_record3_rgb_n_b}) - soc_frame_rgb2ycbcr_yraw);
		soc_frame_rgb2ycbcr_r_minus_yraw <= ($signed({1'd0, soc_frame_rgb2ycbcr_record3_rgb_n_r}) - soc_frame_rgb2ycbcr_yraw);
		soc_frame_rgb2ycbcr_yraw_r0 <= soc_frame_rgb2ycbcr_yraw;
		soc_frame_rgb2ycbcr_cc_mult_ryraw <= (soc_frame_rgb2ycbcr_b_minus_yraw * $signed({1'd0, 8'd141}));
		soc_frame_rgb2ycbcr_cd_mult_byraw <= (soc_frame_rgb2ycbcr_r_minus_yraw * $signed({1'd0, 8'd166}));
		soc_frame_rgb2ycbcr_yraw_r1 <= soc_frame_rgb2ycbcr_yraw_r0;
		soc_frame_rgb2ycbcr_y <= (soc_frame_rgb2ycbcr_yraw_r1 + $signed({1'd0, 5'd16}));
		soc_frame_rgb2ycbcr_cb <= (soc_frame_rgb2ycbcr_cc_mult_ryraw[19:8] + $signed({1'd0, 8'd128}));
		soc_frame_rgb2ycbcr_cr <= (soc_frame_rgb2ycbcr_cd_mult_byraw[19:8] + $signed({1'd0, 8'd128}));
		if ((soc_frame_rgb2ycbcr_y > $signed({1'd0, 8'd255}))) begin
			soc_frame_rgb2ycbcr_source_y <= 8'd255;
		end else begin
			if ((soc_frame_rgb2ycbcr_y < $signed({1'd0, 1'd0}))) begin
				soc_frame_rgb2ycbcr_source_y <= 1'd0;
			end else begin
				soc_frame_rgb2ycbcr_source_y <= soc_frame_rgb2ycbcr_y;
			end
		end
		if ((soc_frame_rgb2ycbcr_cb > $signed({1'd0, 8'd255}))) begin
			soc_frame_rgb2ycbcr_source_cb <= 8'd255;
		end else begin
			if ((soc_frame_rgb2ycbcr_cb < $signed({1'd0, 1'd0}))) begin
				soc_frame_rgb2ycbcr_source_cb <= 1'd0;
			end else begin
				soc_frame_rgb2ycbcr_source_cb <= soc_frame_rgb2ycbcr_cb;
			end
		end
		if ((soc_frame_rgb2ycbcr_cr > $signed({1'd0, 8'd255}))) begin
			soc_frame_rgb2ycbcr_source_cr <= 8'd255;
		end else begin
			if ((soc_frame_rgb2ycbcr_cr < $signed({1'd0, 1'd0}))) begin
				soc_frame_rgb2ycbcr_source_cr <= 1'd0;
			end else begin
				soc_frame_rgb2ycbcr_source_cr <= soc_frame_rgb2ycbcr_cr;
			end
		end
	end
	if (soc_frame_chroma_downsampler_pipe_ce) begin
		soc_frame_chroma_downsampler_valid_n0 <= soc_frame_chroma_downsampler_sink_valid;
	end
	if (soc_frame_chroma_downsampler_pipe_ce) begin
		soc_frame_chroma_downsampler_valid_n1 <= soc_frame_chroma_downsampler_valid_n0;
	end
	if (soc_frame_chroma_downsampler_pipe_ce) begin
		soc_frame_chroma_downsampler_valid_n2 <= soc_frame_chroma_downsampler_valid_n1;
	end
	if (soc_frame_chroma_downsampler_pipe_ce) begin
		soc_frame_chroma_downsampler_first_n0 <= (soc_frame_chroma_downsampler_sink_valid & soc_frame_chroma_downsampler_sink_first);
		soc_frame_chroma_downsampler_last_n0 <= (soc_frame_chroma_downsampler_sink_valid & soc_frame_chroma_downsampler_sink_last);
	end
	if (soc_frame_chroma_downsampler_pipe_ce) begin
		soc_frame_chroma_downsampler_first_n1 <= soc_frame_chroma_downsampler_first_n0;
		soc_frame_chroma_downsampler_last_n1 <= soc_frame_chroma_downsampler_last_n0;
	end
	if (soc_frame_chroma_downsampler_pipe_ce) begin
		soc_frame_chroma_downsampler_first_n2 <= soc_frame_chroma_downsampler_first_n1;
		soc_frame_chroma_downsampler_last_n2 <= soc_frame_chroma_downsampler_last_n1;
	end
	if (soc_frame_chroma_downsampler_ce) begin
		soc_frame_chroma_downsampler_record0_ycbcr_n_y <= soc_frame_chroma_downsampler_sink_y;
		soc_frame_chroma_downsampler_record0_ycbcr_n_cb <= soc_frame_chroma_downsampler_sink_cb;
		soc_frame_chroma_downsampler_record0_ycbcr_n_cr <= soc_frame_chroma_downsampler_sink_cr;
		soc_frame_chroma_downsampler_record1_ycbcr_n_y <= soc_frame_chroma_downsampler_record0_ycbcr_n_y;
		soc_frame_chroma_downsampler_record1_ycbcr_n_cb <= soc_frame_chroma_downsampler_record0_ycbcr_n_cb;
		soc_frame_chroma_downsampler_record1_ycbcr_n_cr <= soc_frame_chroma_downsampler_record0_ycbcr_n_cr;
		soc_frame_chroma_downsampler_record2_ycbcr_n_y <= soc_frame_chroma_downsampler_record1_ycbcr_n_y;
		soc_frame_chroma_downsampler_record2_ycbcr_n_cb <= soc_frame_chroma_downsampler_record1_ycbcr_n_cb;
		soc_frame_chroma_downsampler_record2_ycbcr_n_cr <= soc_frame_chroma_downsampler_record1_ycbcr_n_cr;
		if ((soc_frame_chroma_downsampler_first | (~soc_frame_chroma_downsampler_parity))) begin
			soc_frame_chroma_downsampler_parity <= 1'd1;
		end else begin
			soc_frame_chroma_downsampler_parity <= 1'd0;
		end
		if (soc_frame_chroma_downsampler_parity) begin
			soc_frame_chroma_downsampler_cb_sum <= (soc_frame_chroma_downsampler_sink_cb + soc_frame_chroma_downsampler_record0_ycbcr_n_cb);
			soc_frame_chroma_downsampler_cr_sum <= (soc_frame_chroma_downsampler_sink_cr + soc_frame_chroma_downsampler_record0_ycbcr_n_cr);
		end
		if (soc_frame_chroma_downsampler_parity) begin
			soc_frame_chroma_downsampler_source_y <= soc_frame_chroma_downsampler_record1_ycbcr_n_y;
			soc_frame_chroma_downsampler_source_cb_cr <= soc_frame_chroma_downsampler_cr_mean;
		end else begin
			soc_frame_chroma_downsampler_source_y <= soc_frame_chroma_downsampler_record1_ycbcr_n_y;
			soc_frame_chroma_downsampler_source_cb_cr <= soc_frame_chroma_downsampler_cb_mean;
		end
	end
	soc_frame_fifo_graycounter0_q_binary <= soc_frame_fifo_graycounter0_q_next_binary;
	soc_frame_fifo_graycounter0_q <= soc_frame_fifo_graycounter0_q_next;
	soc_frame_overflow_reset_toggle_o_r <= soc_frame_overflow_reset_toggle_o;
	if (soc_frame_overflow_reset_ack_i) begin
		soc_frame_overflow_reset_ack_toggle_i <= (~soc_frame_overflow_reset_ack_toggle_i);
	end
	if (hdmi_in0_pix_rst) begin
		soc_charsync0_synced <= 1'd0;
		soc_charsync0_data <= 10'd0;
		soc_charsync0_raw_data1 <= 10'd0;
		soc_charsync0_found_control <= 1'd0;
		soc_charsync0_control_position <= 4'd0;
		soc_charsync0_control_counter <= 3'd0;
		soc_charsync0_previous_control_position <= 4'd0;
		soc_charsync0_word_sel <= 4'd0;
		soc_wer0_data_r <= 9'd0;
		soc_wer0_transition_count <= 4'd0;
		soc_wer0_is_control <= 1'd0;
		soc_wer0_is_error <= 1'd0;
		soc_wer0_period_counter <= 24'd0;
		soc_wer0_period_done <= 1'd0;
		soc_wer0_wer_counter <= 24'd0;
		soc_wer0_wer_counter_r <= 24'd0;
		soc_wer0_wer_counter_r_updated <= 1'd0;
		soc_decoding0_valid_o <= 1'd0;
		soc_decoding0_output_d <= 8'd0;
		soc_decoding0_output_c <= 2'd0;
		soc_decoding0_output_de <= 1'd0;
		soc_charsync1_synced <= 1'd0;
		soc_charsync1_data <= 10'd0;
		soc_charsync1_raw_data1 <= 10'd0;
		soc_charsync1_found_control <= 1'd0;
		soc_charsync1_control_position <= 4'd0;
		soc_charsync1_control_counter <= 3'd0;
		soc_charsync1_previous_control_position <= 4'd0;
		soc_charsync1_word_sel <= 4'd0;
		soc_wer1_data_r <= 9'd0;
		soc_wer1_transition_count <= 4'd0;
		soc_wer1_is_control <= 1'd0;
		soc_wer1_is_error <= 1'd0;
		soc_wer1_period_counter <= 24'd0;
		soc_wer1_period_done <= 1'd0;
		soc_wer1_wer_counter <= 24'd0;
		soc_wer1_wer_counter_r <= 24'd0;
		soc_wer1_wer_counter_r_updated <= 1'd0;
		soc_decoding1_valid_o <= 1'd0;
		soc_decoding1_output_d <= 8'd0;
		soc_decoding1_output_c <= 2'd0;
		soc_decoding1_output_de <= 1'd0;
		soc_charsync2_synced <= 1'd0;
		soc_charsync2_data <= 10'd0;
		soc_charsync2_raw_data1 <= 10'd0;
		soc_charsync2_found_control <= 1'd0;
		soc_charsync2_control_position <= 4'd0;
		soc_charsync2_control_counter <= 3'd0;
		soc_charsync2_previous_control_position <= 4'd0;
		soc_charsync2_word_sel <= 4'd0;
		soc_wer2_data_r <= 9'd0;
		soc_wer2_transition_count <= 4'd0;
		soc_wer2_is_control <= 1'd0;
		soc_wer2_is_error <= 1'd0;
		soc_wer2_period_counter <= 24'd0;
		soc_wer2_period_done <= 1'd0;
		soc_wer2_wer_counter <= 24'd0;
		soc_wer2_wer_counter_r <= 24'd0;
		soc_wer2_wer_counter_r_updated <= 1'd0;
		soc_decoding2_valid_o <= 1'd0;
		soc_decoding2_output_d <= 8'd0;
		soc_decoding2_output_c <= 2'd0;
		soc_decoding2_output_de <= 1'd0;
		soc_chansync_chan_synced <= 1'd0;
		soc_chansync_syncbuffer0_produce <= 3'd0;
		soc_chansync_syncbuffer0_consume <= 3'd0;
		soc_chansync_syncbuffer1_produce <= 3'd0;
		soc_chansync_syncbuffer1_consume <= 3'd0;
		soc_chansync_syncbuffer2_produce <= 3'd0;
		soc_chansync_syncbuffer2_consume <= 3'd0;
		soc_syncpol_valid_o <= 1'd0;
		soc_syncpol_r <= 8'd0;
		soc_syncpol_g <= 8'd0;
		soc_syncpol_b <= 8'd0;
		soc_syncpol_de_r <= 1'd0;
		soc_syncpol_c_polarity <= 2'd0;
		soc_syncpol_c_out <= 2'd0;
		soc_resdetection_de_r <= 1'd0;
		soc_resdetection_hcounter <= 11'd0;
		soc_resdetection_hcounter_st <= 11'd0;
		soc_resdetection_vsync_r <= 1'd0;
		soc_resdetection_vcounter <= 11'd0;
		soc_resdetection_vcounter_st <= 11'd0;
		soc_frame_de_r <= 1'd0;
		soc_frame_rgb2ycbcr_source_y <= 8'd0;
		soc_frame_rgb2ycbcr_source_cb <= 8'd0;
		soc_frame_rgb2ycbcr_source_cr <= 8'd0;
		soc_frame_rgb2ycbcr_record0_rgb_n_r <= 8'd0;
		soc_frame_rgb2ycbcr_record0_rgb_n_g <= 8'd0;
		soc_frame_rgb2ycbcr_record0_rgb_n_b <= 8'd0;
		soc_frame_rgb2ycbcr_record1_rgb_n_r <= 8'd0;
		soc_frame_rgb2ycbcr_record1_rgb_n_g <= 8'd0;
		soc_frame_rgb2ycbcr_record1_rgb_n_b <= 8'd0;
		soc_frame_rgb2ycbcr_record2_rgb_n_r <= 8'd0;
		soc_frame_rgb2ycbcr_record2_rgb_n_g <= 8'd0;
		soc_frame_rgb2ycbcr_record2_rgb_n_b <= 8'd0;
		soc_frame_rgb2ycbcr_record3_rgb_n_r <= 8'd0;
		soc_frame_rgb2ycbcr_record3_rgb_n_g <= 8'd0;
		soc_frame_rgb2ycbcr_record3_rgb_n_b <= 8'd0;
		soc_frame_rgb2ycbcr_record4_rgb_n_r <= 8'd0;
		soc_frame_rgb2ycbcr_record4_rgb_n_g <= 8'd0;
		soc_frame_rgb2ycbcr_record4_rgb_n_b <= 8'd0;
		soc_frame_rgb2ycbcr_record5_rgb_n_r <= 8'd0;
		soc_frame_rgb2ycbcr_record5_rgb_n_g <= 8'd0;
		soc_frame_rgb2ycbcr_record5_rgb_n_b <= 8'd0;
		soc_frame_rgb2ycbcr_record6_rgb_n_r <= 8'd0;
		soc_frame_rgb2ycbcr_record6_rgb_n_g <= 8'd0;
		soc_frame_rgb2ycbcr_record6_rgb_n_b <= 8'd0;
		soc_frame_rgb2ycbcr_record7_rgb_n_r <= 8'd0;
		soc_frame_rgb2ycbcr_record7_rgb_n_g <= 8'd0;
		soc_frame_rgb2ycbcr_record7_rgb_n_b <= 8'd0;
		soc_frame_rgb2ycbcr_r_minus_g <= 9'sd512;
		soc_frame_rgb2ycbcr_b_minus_g <= 9'sd512;
		soc_frame_rgb2ycbcr_ca_mult_rg <= 17'sd131072;
		soc_frame_rgb2ycbcr_cb_mult_bg <= 17'sd131072;
		soc_frame_rgb2ycbcr_carg_plus_cbbg <= 25'sd33554432;
		soc_frame_rgb2ycbcr_yraw <= 11'sd2048;
		soc_frame_rgb2ycbcr_b_minus_yraw <= 12'sd4096;
		soc_frame_rgb2ycbcr_r_minus_yraw <= 12'sd4096;
		soc_frame_rgb2ycbcr_yraw_r0 <= 11'sd2048;
		soc_frame_rgb2ycbcr_cc_mult_ryraw <= 20'sd1048576;
		soc_frame_rgb2ycbcr_cd_mult_byraw <= 20'sd1048576;
		soc_frame_rgb2ycbcr_yraw_r1 <= 11'sd2048;
		soc_frame_rgb2ycbcr_y <= 11'sd2048;
		soc_frame_rgb2ycbcr_cb <= 12'sd4096;
		soc_frame_rgb2ycbcr_cr <= 12'sd4096;
		soc_frame_rgb2ycbcr_valid_n0 <= 1'd0;
		soc_frame_rgb2ycbcr_valid_n1 <= 1'd0;
		soc_frame_rgb2ycbcr_valid_n2 <= 1'd0;
		soc_frame_rgb2ycbcr_valid_n3 <= 1'd0;
		soc_frame_rgb2ycbcr_valid_n4 <= 1'd0;
		soc_frame_rgb2ycbcr_valid_n5 <= 1'd0;
		soc_frame_rgb2ycbcr_valid_n6 <= 1'd0;
		soc_frame_rgb2ycbcr_valid_n7 <= 1'd0;
		soc_frame_rgb2ycbcr_first_n0 <= 1'd0;
		soc_frame_rgb2ycbcr_last_n0 <= 1'd0;
		soc_frame_rgb2ycbcr_first_n1 <= 1'd0;
		soc_frame_rgb2ycbcr_last_n1 <= 1'd0;
		soc_frame_rgb2ycbcr_first_n2 <= 1'd0;
		soc_frame_rgb2ycbcr_last_n2 <= 1'd0;
		soc_frame_rgb2ycbcr_first_n3 <= 1'd0;
		soc_frame_rgb2ycbcr_last_n3 <= 1'd0;
		soc_frame_rgb2ycbcr_first_n4 <= 1'd0;
		soc_frame_rgb2ycbcr_last_n4 <= 1'd0;
		soc_frame_rgb2ycbcr_first_n5 <= 1'd0;
		soc_frame_rgb2ycbcr_last_n5 <= 1'd0;
		soc_frame_rgb2ycbcr_first_n6 <= 1'd0;
		soc_frame_rgb2ycbcr_last_n6 <= 1'd0;
		soc_frame_rgb2ycbcr_first_n7 <= 1'd0;
		soc_frame_rgb2ycbcr_last_n7 <= 1'd0;
		soc_frame_chroma_downsampler_source_y <= 8'd0;
		soc_frame_chroma_downsampler_source_cb_cr <= 8'd0;
		soc_frame_chroma_downsampler_record0_ycbcr_n_y <= 8'd0;
		soc_frame_chroma_downsampler_record0_ycbcr_n_cb <= 8'd0;
		soc_frame_chroma_downsampler_record0_ycbcr_n_cr <= 8'd0;
		soc_frame_chroma_downsampler_record1_ycbcr_n_y <= 8'd0;
		soc_frame_chroma_downsampler_record1_ycbcr_n_cb <= 8'd0;
		soc_frame_chroma_downsampler_record1_ycbcr_n_cr <= 8'd0;
		soc_frame_chroma_downsampler_record2_ycbcr_n_y <= 8'd0;
		soc_frame_chroma_downsampler_record2_ycbcr_n_cb <= 8'd0;
		soc_frame_chroma_downsampler_record2_ycbcr_n_cr <= 8'd0;
		soc_frame_chroma_downsampler_parity <= 1'd0;
		soc_frame_chroma_downsampler_cb_sum <= 9'd0;
		soc_frame_chroma_downsampler_cr_sum <= 9'd0;
		soc_frame_chroma_downsampler_valid_n0 <= 1'd0;
		soc_frame_chroma_downsampler_valid_n1 <= 1'd0;
		soc_frame_chroma_downsampler_valid_n2 <= 1'd0;
		soc_frame_chroma_downsampler_first_n0 <= 1'd0;
		soc_frame_chroma_downsampler_last_n0 <= 1'd0;
		soc_frame_chroma_downsampler_first_n1 <= 1'd0;
		soc_frame_chroma_downsampler_last_n1 <= 1'd0;
		soc_frame_chroma_downsampler_first_n2 <= 1'd0;
		soc_frame_chroma_downsampler_last_n2 <= 1'd0;
		soc_frame_next_de0 <= 1'd0;
		soc_frame_next_vsync0 <= 1'd0;
		soc_frame_next_de1 <= 1'd0;
		soc_frame_next_vsync1 <= 1'd0;
		soc_frame_next_de2 <= 1'd0;
		soc_frame_next_vsync2 <= 1'd0;
		soc_frame_next_de3 <= 1'd0;
		soc_frame_next_vsync3 <= 1'd0;
		soc_frame_next_de4 <= 1'd0;
		soc_frame_next_vsync4 <= 1'd0;
		soc_frame_next_de5 <= 1'd0;
		soc_frame_next_vsync5 <= 1'd0;
		soc_frame_next_de6 <= 1'd0;
		soc_frame_next_vsync6 <= 1'd0;
		soc_frame_next_de7 <= 1'd0;
		soc_frame_next_vsync7 <= 1'd0;
		soc_frame_next_de8 <= 1'd0;
		soc_frame_next_vsync8 <= 1'd0;
		soc_frame_next_de9 <= 1'd0;
		soc_frame_next_vsync9 <= 1'd0;
		soc_frame_next_de10 <= 1'd0;
		soc_frame_next_vsync10 <= 1'd0;
		soc_frame_vsync_r <= 1'd0;
		soc_frame_cur_word <= 128'd0;
		soc_frame_cur_word_valid <= 1'd0;
		soc_frame_pack_counter <= 3'd0;
		soc_frame_fifo_graycounter0_q <= 10'd0;
		soc_frame_fifo_graycounter0_q_binary <= 10'd0;
		soc_frame_pix_overflow <= 1'd0;
	end
	vns_xilinxmultiregimpl43_regs0 <= soc_frame_fifo_graycounter1_q;
	vns_xilinxmultiregimpl43_regs1 <= vns_xilinxmultiregimpl43_regs0;
	vns_xilinxmultiregimpl45_regs0 <= soc_frame_overflow_reset_toggle_i;
	vns_xilinxmultiregimpl45_regs1 <= vns_xilinxmultiregimpl45_regs0;
end

always @(posedge hdmi_out0_pix_clk) begin
	soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_binary <= soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next_binary;
	soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q <= soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_next;
	soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_binary <= soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next_binary;
	soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q <= soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_next;
	if (soc_hdmi_out0_dram_port_counter_ce) begin
		soc_hdmi_out0_dram_port_counter <= (soc_hdmi_out0_dram_port_counter + 1'd1);
	end
	if ((soc_hdmi_out0_dram_port_rdata_converter_source_valid & soc_hdmi_out0_dram_port_rdata_converter_source_ready)) begin
		soc_hdmi_out0_dram_port_rdata_chunk <= {soc_hdmi_out0_dram_port_rdata_chunk[6:0], soc_hdmi_out0_dram_port_rdata_chunk[7]};
	end
	if (((soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_we & soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_writable) & (~soc_hdmi_out0_dram_port_cmd_buffer_replace))) begin
		soc_hdmi_out0_dram_port_cmd_buffer_produce <= (soc_hdmi_out0_dram_port_cmd_buffer_produce + 1'd1);
	end
	if (soc_hdmi_out0_dram_port_cmd_buffer_do_read) begin
		soc_hdmi_out0_dram_port_cmd_buffer_consume <= (soc_hdmi_out0_dram_port_cmd_buffer_consume + 1'd1);
	end
	if (((soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_we & soc_hdmi_out0_dram_port_cmd_buffer_syncfifo_writable) & (~soc_hdmi_out0_dram_port_cmd_buffer_replace))) begin
		if ((~soc_hdmi_out0_dram_port_cmd_buffer_do_read)) begin
			soc_hdmi_out0_dram_port_cmd_buffer_level <= (soc_hdmi_out0_dram_port_cmd_buffer_level + 1'd1);
		end
	end else begin
		if (soc_hdmi_out0_dram_port_cmd_buffer_do_read) begin
			soc_hdmi_out0_dram_port_cmd_buffer_level <= (soc_hdmi_out0_dram_port_cmd_buffer_level - 1'd1);
		end
	end
	if (soc_hdmi_out0_dram_port_rdata_buffer_pipe_ce) begin
		soc_hdmi_out0_dram_port_rdata_buffer_valid_n <= soc_hdmi_out0_dram_port_rdata_buffer_sink_valid;
	end
	if (soc_hdmi_out0_dram_port_rdata_buffer_pipe_ce) begin
		soc_hdmi_out0_dram_port_rdata_buffer_first_n <= (soc_hdmi_out0_dram_port_rdata_buffer_sink_valid & soc_hdmi_out0_dram_port_rdata_buffer_sink_first);
		soc_hdmi_out0_dram_port_rdata_buffer_last_n <= (soc_hdmi_out0_dram_port_rdata_buffer_sink_valid & soc_hdmi_out0_dram_port_rdata_buffer_sink_last);
	end
	if (soc_hdmi_out0_dram_port_rdata_buffer_pipe_ce) begin
		soc_hdmi_out0_dram_port_rdata_buffer_source_payload_data <= soc_hdmi_out0_dram_port_rdata_buffer_sink_payload_data;
	end
	if ((soc_hdmi_out0_dram_port_rdata_converter_converter_source_valid & soc_hdmi_out0_dram_port_rdata_converter_converter_source_ready)) begin
		if (soc_hdmi_out0_dram_port_rdata_converter_converter_last) begin
			soc_hdmi_out0_dram_port_rdata_converter_converter_mux <= 1'd0;
		end else begin
			soc_hdmi_out0_dram_port_rdata_converter_converter_mux <= (soc_hdmi_out0_dram_port_rdata_converter_converter_mux + 1'd1);
		end
	end
	soc_hdmi_out0_de_r <= soc_hdmi_out0_core_source_source_param_de;
	soc_hdmi_out0_core_source_valid_d <= soc_hdmi_out0_core_source_source_valid;
	soc_hdmi_out0_core_source_data_d <= soc_hdmi_out0_core_source_source_payload_data;
	if (soc_hdmi_out0_core_underflow_enable) begin
		if ((~soc_hdmi_out0_core_source_source_valid)) begin
			soc_hdmi_out0_core_underflow_counter <= (soc_hdmi_out0_core_underflow_counter + 1'd1);
		end
	end else begin
		soc_hdmi_out0_core_underflow_counter <= 1'd0;
	end
	if (soc_hdmi_out0_core_underflow_update) begin
		soc_hdmi_out0_core_underflow_counter_status <= soc_hdmi_out0_core_underflow_counter;
	end
	soc_hdmi_out0_core_initiator_cdc_graycounter1_q_binary <= soc_hdmi_out0_core_initiator_cdc_graycounter1_q_next_binary;
	soc_hdmi_out0_core_initiator_cdc_graycounter1_q <= soc_hdmi_out0_core_initiator_cdc_graycounter1_q_next;
	if ((~soc_hdmi_out0_core_timinggenerator_sink_valid)) begin
		soc_hdmi_out0_core_timinggenerator_hactive <= 1'd0;
		soc_hdmi_out0_core_timinggenerator_vactive <= 1'd0;
		soc_hdmi_out0_core_timinggenerator_hcounter <= 1'd0;
		soc_hdmi_out0_core_timinggenerator_vcounter <= 1'd0;
	end else begin
		if (soc_hdmi_out0_core_timinggenerator_source_ready) begin
			soc_hdmi_out0_core_timinggenerator_source_last <= 1'd0;
			soc_hdmi_out0_core_timinggenerator_hcounter <= (soc_hdmi_out0_core_timinggenerator_hcounter + 1'd1);
			if ((soc_hdmi_out0_core_timinggenerator_hcounter == 1'd0)) begin
				soc_hdmi_out0_core_timinggenerator_hactive <= 1'd1;
			end
			if ((soc_hdmi_out0_core_timinggenerator_hcounter == soc_hdmi_out0_core_timinggenerator_sink_payload_hres)) begin
				soc_hdmi_out0_core_timinggenerator_hactive <= 1'd0;
			end
			if ((soc_hdmi_out0_core_timinggenerator_hcounter == soc_hdmi_out0_core_timinggenerator_sink_payload_hsync_start)) begin
				soc_hdmi_out0_core_timinggenerator_source_payload_hsync <= 1'd1;
			end
			if ((soc_hdmi_out0_core_timinggenerator_hcounter == soc_hdmi_out0_core_timinggenerator_sink_payload_hsync_end)) begin
				soc_hdmi_out0_core_timinggenerator_source_payload_hsync <= 1'd0;
			end
			if ((soc_hdmi_out0_core_timinggenerator_hcounter == soc_hdmi_out0_core_timinggenerator_sink_payload_hscan)) begin
				soc_hdmi_out0_core_timinggenerator_hcounter <= 1'd0;
				if ((soc_hdmi_out0_core_timinggenerator_vcounter == soc_hdmi_out0_core_timinggenerator_sink_payload_vscan)) begin
					soc_hdmi_out0_core_timinggenerator_vcounter <= 1'd0;
					soc_hdmi_out0_core_timinggenerator_source_last <= 1'd1;
				end else begin
					soc_hdmi_out0_core_timinggenerator_vcounter <= (soc_hdmi_out0_core_timinggenerator_vcounter + 1'd1);
				end
			end
			if ((soc_hdmi_out0_core_timinggenerator_vcounter == 1'd0)) begin
				soc_hdmi_out0_core_timinggenerator_vactive <= 1'd1;
			end
			if ((soc_hdmi_out0_core_timinggenerator_vcounter == soc_hdmi_out0_core_timinggenerator_sink_payload_vres)) begin
				soc_hdmi_out0_core_timinggenerator_vactive <= 1'd0;
			end
			if ((soc_hdmi_out0_core_timinggenerator_vcounter == soc_hdmi_out0_core_timinggenerator_sink_payload_vsync_start)) begin
				soc_hdmi_out0_core_timinggenerator_source_payload_vsync <= 1'd1;
			end
			if ((soc_hdmi_out0_core_timinggenerator_vcounter == soc_hdmi_out0_core_timinggenerator_sink_payload_vsync_end)) begin
				soc_hdmi_out0_core_timinggenerator_source_payload_vsync <= 1'd0;
			end
		end
	end
	if (soc_hdmi_out0_core_dmareader_request_issued) begin
		if ((~soc_hdmi_out0_core_dmareader_data_dequeued)) begin
			soc_hdmi_out0_core_dmareader_rsv_level <= (soc_hdmi_out0_core_dmareader_rsv_level + 1'd1);
		end
	end else begin
		if (soc_hdmi_out0_core_dmareader_data_dequeued) begin
			soc_hdmi_out0_core_dmareader_rsv_level <= (soc_hdmi_out0_core_dmareader_rsv_level - 1'd1);
		end
	end
	if (soc_hdmi_out0_core_dmareader_fifo_syncfifo_re) begin
		soc_hdmi_out0_core_dmareader_fifo_readable <= 1'd1;
	end else begin
		if (soc_hdmi_out0_core_dmareader_fifo_re) begin
			soc_hdmi_out0_core_dmareader_fifo_readable <= 1'd0;
		end
	end
	if (((soc_hdmi_out0_core_dmareader_fifo_syncfifo_we & soc_hdmi_out0_core_dmareader_fifo_syncfifo_writable) & (~soc_hdmi_out0_core_dmareader_fifo_replace))) begin
		soc_hdmi_out0_core_dmareader_fifo_produce <= (soc_hdmi_out0_core_dmareader_fifo_produce + 1'd1);
	end
	if (soc_hdmi_out0_core_dmareader_fifo_do_read) begin
		soc_hdmi_out0_core_dmareader_fifo_consume <= (soc_hdmi_out0_core_dmareader_fifo_consume + 1'd1);
	end
	if (((soc_hdmi_out0_core_dmareader_fifo_syncfifo_we & soc_hdmi_out0_core_dmareader_fifo_syncfifo_writable) & (~soc_hdmi_out0_core_dmareader_fifo_replace))) begin
		if ((~soc_hdmi_out0_core_dmareader_fifo_do_read)) begin
			soc_hdmi_out0_core_dmareader_fifo_level0 <= (soc_hdmi_out0_core_dmareader_fifo_level0 + 1'd1);
		end
	end else begin
		if (soc_hdmi_out0_core_dmareader_fifo_do_read) begin
			soc_hdmi_out0_core_dmareader_fifo_level0 <= (soc_hdmi_out0_core_dmareader_fifo_level0 - 1'd1);
		end
	end
	vns_videoout_state <= vns_videoout_next_state;
	if (soc_hdmi_out0_core_dmareader_offset_next_value_ce) begin
		soc_hdmi_out0_core_dmareader_offset <= soc_hdmi_out0_core_dmareader_offset_next_value;
	end
	soc_hdmi_out0_core_toggle_o_r <= soc_hdmi_out0_core_toggle_o;
	if ((soc_hdmi_out0_resetinserter_sink_sink_valid & soc_hdmi_out0_resetinserter_sink_sink_ready)) begin
		soc_hdmi_out0_resetinserter_parity_in <= (~soc_hdmi_out0_resetinserter_parity_in);
	end
	if ((soc_hdmi_out0_resetinserter_source_source_valid & soc_hdmi_out0_resetinserter_source_source_ready)) begin
		soc_hdmi_out0_resetinserter_parity_out <= (~soc_hdmi_out0_resetinserter_parity_out);
	end
	if (((soc_hdmi_out0_resetinserter_y_fifo_syncfifo_we & soc_hdmi_out0_resetinserter_y_fifo_syncfifo_writable) & (~soc_hdmi_out0_resetinserter_y_fifo_replace))) begin
		soc_hdmi_out0_resetinserter_y_fifo_produce <= (soc_hdmi_out0_resetinserter_y_fifo_produce + 1'd1);
	end
	if (soc_hdmi_out0_resetinserter_y_fifo_do_read) begin
		soc_hdmi_out0_resetinserter_y_fifo_consume <= (soc_hdmi_out0_resetinserter_y_fifo_consume + 1'd1);
	end
	if (((soc_hdmi_out0_resetinserter_y_fifo_syncfifo_we & soc_hdmi_out0_resetinserter_y_fifo_syncfifo_writable) & (~soc_hdmi_out0_resetinserter_y_fifo_replace))) begin
		if ((~soc_hdmi_out0_resetinserter_y_fifo_do_read)) begin
			soc_hdmi_out0_resetinserter_y_fifo_level <= (soc_hdmi_out0_resetinserter_y_fifo_level + 1'd1);
		end
	end else begin
		if (soc_hdmi_out0_resetinserter_y_fifo_do_read) begin
			soc_hdmi_out0_resetinserter_y_fifo_level <= (soc_hdmi_out0_resetinserter_y_fifo_level - 1'd1);
		end
	end
	if (((soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_we & soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_writable) & (~soc_hdmi_out0_resetinserter_cb_fifo_replace))) begin
		soc_hdmi_out0_resetinserter_cb_fifo_produce <= (soc_hdmi_out0_resetinserter_cb_fifo_produce + 1'd1);
	end
	if (soc_hdmi_out0_resetinserter_cb_fifo_do_read) begin
		soc_hdmi_out0_resetinserter_cb_fifo_consume <= (soc_hdmi_out0_resetinserter_cb_fifo_consume + 1'd1);
	end
	if (((soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_we & soc_hdmi_out0_resetinserter_cb_fifo_syncfifo_writable) & (~soc_hdmi_out0_resetinserter_cb_fifo_replace))) begin
		if ((~soc_hdmi_out0_resetinserter_cb_fifo_do_read)) begin
			soc_hdmi_out0_resetinserter_cb_fifo_level <= (soc_hdmi_out0_resetinserter_cb_fifo_level + 1'd1);
		end
	end else begin
		if (soc_hdmi_out0_resetinserter_cb_fifo_do_read) begin
			soc_hdmi_out0_resetinserter_cb_fifo_level <= (soc_hdmi_out0_resetinserter_cb_fifo_level - 1'd1);
		end
	end
	if (((soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_we & soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_writable) & (~soc_hdmi_out0_resetinserter_cr_fifo_replace))) begin
		soc_hdmi_out0_resetinserter_cr_fifo_produce <= (soc_hdmi_out0_resetinserter_cr_fifo_produce + 1'd1);
	end
	if (soc_hdmi_out0_resetinserter_cr_fifo_do_read) begin
		soc_hdmi_out0_resetinserter_cr_fifo_consume <= (soc_hdmi_out0_resetinserter_cr_fifo_consume + 1'd1);
	end
	if (((soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_we & soc_hdmi_out0_resetinserter_cr_fifo_syncfifo_writable) & (~soc_hdmi_out0_resetinserter_cr_fifo_replace))) begin
		if ((~soc_hdmi_out0_resetinserter_cr_fifo_do_read)) begin
			soc_hdmi_out0_resetinserter_cr_fifo_level <= (soc_hdmi_out0_resetinserter_cr_fifo_level + 1'd1);
		end
	end else begin
		if (soc_hdmi_out0_resetinserter_cr_fifo_do_read) begin
			soc_hdmi_out0_resetinserter_cr_fifo_level <= (soc_hdmi_out0_resetinserter_cr_fifo_level - 1'd1);
		end
	end
	if (soc_hdmi_out0_resetinserter_reset) begin
		soc_hdmi_out0_resetinserter_y_fifo_level <= 3'd0;
		soc_hdmi_out0_resetinserter_y_fifo_produce <= 2'd0;
		soc_hdmi_out0_resetinserter_y_fifo_consume <= 2'd0;
		soc_hdmi_out0_resetinserter_cb_fifo_level <= 3'd0;
		soc_hdmi_out0_resetinserter_cb_fifo_produce <= 2'd0;
		soc_hdmi_out0_resetinserter_cb_fifo_consume <= 2'd0;
		soc_hdmi_out0_resetinserter_cr_fifo_level <= 3'd0;
		soc_hdmi_out0_resetinserter_cr_fifo_produce <= 2'd0;
		soc_hdmi_out0_resetinserter_cr_fifo_consume <= 2'd0;
		soc_hdmi_out0_resetinserter_parity_in <= 1'd0;
		soc_hdmi_out0_resetinserter_parity_out <= 1'd0;
	end
	if (soc_hdmi_out0_pipe_ce) begin
		soc_hdmi_out0_valid_n0 <= soc_hdmi_out0_sink_valid;
	end
	if (soc_hdmi_out0_pipe_ce) begin
		soc_hdmi_out0_valid_n1 <= soc_hdmi_out0_valid_n0;
	end
	if (soc_hdmi_out0_pipe_ce) begin
		soc_hdmi_out0_valid_n2 <= soc_hdmi_out0_valid_n1;
	end
	if (soc_hdmi_out0_pipe_ce) begin
		soc_hdmi_out0_valid_n3 <= soc_hdmi_out0_valid_n2;
	end
	if (soc_hdmi_out0_pipe_ce) begin
		soc_hdmi_out0_first_n0 <= (soc_hdmi_out0_sink_valid & soc_hdmi_out0_sink_first);
		soc_hdmi_out0_last_n0 <= (soc_hdmi_out0_sink_valid & soc_hdmi_out0_sink_last);
	end
	if (soc_hdmi_out0_pipe_ce) begin
		soc_hdmi_out0_first_n1 <= soc_hdmi_out0_first_n0;
		soc_hdmi_out0_last_n1 <= soc_hdmi_out0_last_n0;
	end
	if (soc_hdmi_out0_pipe_ce) begin
		soc_hdmi_out0_first_n2 <= soc_hdmi_out0_first_n1;
		soc_hdmi_out0_last_n2 <= soc_hdmi_out0_last_n1;
	end
	if (soc_hdmi_out0_pipe_ce) begin
		soc_hdmi_out0_first_n3 <= soc_hdmi_out0_first_n2;
		soc_hdmi_out0_last_n3 <= soc_hdmi_out0_last_n2;
	end
	if (soc_hdmi_out0_ce) begin
		soc_hdmi_out0_record0_ycbcr_n_y <= soc_hdmi_out0_sink_y;
		soc_hdmi_out0_record0_ycbcr_n_cb <= soc_hdmi_out0_sink_cb;
		soc_hdmi_out0_record0_ycbcr_n_cr <= soc_hdmi_out0_sink_cr;
		soc_hdmi_out0_record1_ycbcr_n_y <= soc_hdmi_out0_record0_ycbcr_n_y;
		soc_hdmi_out0_record1_ycbcr_n_cb <= soc_hdmi_out0_record0_ycbcr_n_cb;
		soc_hdmi_out0_record1_ycbcr_n_cr <= soc_hdmi_out0_record0_ycbcr_n_cr;
		soc_hdmi_out0_record2_ycbcr_n_y <= soc_hdmi_out0_record1_ycbcr_n_y;
		soc_hdmi_out0_record2_ycbcr_n_cb <= soc_hdmi_out0_record1_ycbcr_n_cb;
		soc_hdmi_out0_record2_ycbcr_n_cr <= soc_hdmi_out0_record1_ycbcr_n_cr;
		soc_hdmi_out0_record3_ycbcr_n_y <= soc_hdmi_out0_record2_ycbcr_n_y;
		soc_hdmi_out0_record3_ycbcr_n_cb <= soc_hdmi_out0_record2_ycbcr_n_cb;
		soc_hdmi_out0_record3_ycbcr_n_cr <= soc_hdmi_out0_record2_ycbcr_n_cr;
		soc_hdmi_out0_cb_minus_coffset <= (soc_hdmi_out0_sink_cb - 8'd128);
		soc_hdmi_out0_cr_minus_coffset <= (soc_hdmi_out0_sink_cr - 8'd128);
		soc_hdmi_out0_y_minus_yoffset <= (soc_hdmi_out0_record0_ycbcr_n_y - 5'd16);
		soc_hdmi_out0_cr_minus_coffset_mult_acoef <= (soc_hdmi_out0_cr_minus_coffset * $signed({1'd0, 7'd98}));
		soc_hdmi_out0_cb_minus_coffset_mult_bcoef <= (soc_hdmi_out0_cb_minus_coffset * 5'sd23);
		soc_hdmi_out0_cr_minus_coffset_mult_ccoef <= (soc_hdmi_out0_cr_minus_coffset * 6'sd41);
		soc_hdmi_out0_cb_minus_coffset_mult_dcoef <= (soc_hdmi_out0_cb_minus_coffset * $signed({1'd0, 7'd116}));
		soc_hdmi_out0_r <= (soc_hdmi_out0_y_minus_yoffset + soc_hdmi_out0_cr_minus_coffset_mult_acoef[19:6]);
		soc_hdmi_out0_g <= ((soc_hdmi_out0_y_minus_yoffset + soc_hdmi_out0_cb_minus_coffset_mult_bcoef[19:6]) + soc_hdmi_out0_cr_minus_coffset_mult_ccoef[19:6]);
		soc_hdmi_out0_b <= (soc_hdmi_out0_y_minus_yoffset + soc_hdmi_out0_cb_minus_coffset_mult_dcoef[19:6]);
		if ((soc_hdmi_out0_r > $signed({1'd0, 8'd255}))) begin
			soc_hdmi_out0_source_r <= 8'd255;
		end else begin
			if ((soc_hdmi_out0_r < $signed({1'd0, 1'd0}))) begin
				soc_hdmi_out0_source_r <= 1'd0;
			end else begin
				soc_hdmi_out0_source_r <= soc_hdmi_out0_r;
			end
		end
		if ((soc_hdmi_out0_g > $signed({1'd0, 8'd255}))) begin
			soc_hdmi_out0_source_g <= 8'd255;
		end else begin
			if ((soc_hdmi_out0_g < $signed({1'd0, 1'd0}))) begin
				soc_hdmi_out0_source_g <= 1'd0;
			end else begin
				soc_hdmi_out0_source_g <= soc_hdmi_out0_g;
			end
		end
		if ((soc_hdmi_out0_b > $signed({1'd0, 8'd255}))) begin
			soc_hdmi_out0_source_b <= 8'd255;
		end else begin
			if ((soc_hdmi_out0_b < $signed({1'd0, 1'd0}))) begin
				soc_hdmi_out0_source_b <= 1'd0;
			end else begin
				soc_hdmi_out0_source_b <= soc_hdmi_out0_b;
			end
		end
	end
	soc_hdmi_out0_next_s0 <= soc_hdmi_out0_sink_payload_hsync;
	soc_hdmi_out0_next_s1 <= soc_hdmi_out0_next_s0;
	soc_hdmi_out0_next_s2 <= soc_hdmi_out0_next_s1;
	soc_hdmi_out0_next_s3 <= soc_hdmi_out0_next_s2;
	soc_hdmi_out0_next_s4 <= soc_hdmi_out0_next_s3;
	soc_hdmi_out0_next_s5 <= soc_hdmi_out0_next_s4;
	soc_hdmi_out0_next_s6 <= soc_hdmi_out0_sink_payload_vsync;
	soc_hdmi_out0_next_s7 <= soc_hdmi_out0_next_s6;
	soc_hdmi_out0_next_s8 <= soc_hdmi_out0_next_s7;
	soc_hdmi_out0_next_s9 <= soc_hdmi_out0_next_s8;
	soc_hdmi_out0_next_s10 <= soc_hdmi_out0_next_s9;
	soc_hdmi_out0_next_s11 <= soc_hdmi_out0_next_s10;
	soc_hdmi_out0_next_s12 <= soc_hdmi_out0_sink_payload_de;
	soc_hdmi_out0_next_s13 <= soc_hdmi_out0_next_s12;
	soc_hdmi_out0_next_s14 <= soc_hdmi_out0_next_s13;
	soc_hdmi_out0_next_s15 <= soc_hdmi_out0_next_s14;
	soc_hdmi_out0_next_s16 <= soc_hdmi_out0_next_s15;
	soc_hdmi_out0_next_s17 <= soc_hdmi_out0_next_s16;
	soc_hdmi_out0_driver_s7hdmioutclocking_ce <= (~hdmi_out0_pix_rst);
	soc_hdmi_out0_driver_hdmi_phy_es0_ce <= (~hdmi_out0_pix_rst);
	soc_hdmi_out0_driver_hdmi_phy_es0_n1d <= (((((((soc_hdmi_out0_driver_hdmi_phy_es0_d0[0] + soc_hdmi_out0_driver_hdmi_phy_es0_d0[1]) + soc_hdmi_out0_driver_hdmi_phy_es0_d0[2]) + soc_hdmi_out0_driver_hdmi_phy_es0_d0[3]) + soc_hdmi_out0_driver_hdmi_phy_es0_d0[4]) + soc_hdmi_out0_driver_hdmi_phy_es0_d0[5]) + soc_hdmi_out0_driver_hdmi_phy_es0_d0[6]) + soc_hdmi_out0_driver_hdmi_phy_es0_d0[7]);
	soc_hdmi_out0_driver_hdmi_phy_es0_d1 <= soc_hdmi_out0_driver_hdmi_phy_es0_d0;
	soc_hdmi_out0_driver_hdmi_phy_es0_q_m[0] <= soc_hdmi_out0_driver_hdmi_phy_es0_d1[0];
	soc_hdmi_out0_driver_hdmi_phy_es0_q_m[1] <= ((soc_hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es0_q_m[2] <= ((((soc_hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es0_q_m[3] <= ((((((soc_hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[3]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es0_q_m[4] <= ((((((((soc_hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[3]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[4]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es0_q_m[5] <= ((((((((((soc_hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[3]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[4]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[5]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es0_q_m[6] <= ((((((((((((soc_hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[3]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[4]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[5]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[6]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es0_q_m[7] <= ((((((((((((((soc_hdmi_out0_driver_hdmi_phy_es0_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[3]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[4]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[5]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[6]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es0_d1[7]) ^ soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es0_q_m[8] <= (~soc_hdmi_out0_driver_hdmi_phy_es0_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es0_n0q_m <= ((((((((~soc_hdmi_out0_driver_hdmi_phy_es0_q_m[0]) + (~soc_hdmi_out0_driver_hdmi_phy_es0_q_m[1])) + (~soc_hdmi_out0_driver_hdmi_phy_es0_q_m[2])) + (~soc_hdmi_out0_driver_hdmi_phy_es0_q_m[3])) + (~soc_hdmi_out0_driver_hdmi_phy_es0_q_m[4])) + (~soc_hdmi_out0_driver_hdmi_phy_es0_q_m[5])) + (~soc_hdmi_out0_driver_hdmi_phy_es0_q_m[6])) + (~soc_hdmi_out0_driver_hdmi_phy_es0_q_m[7]));
	soc_hdmi_out0_driver_hdmi_phy_es0_n1q_m <= (((((((soc_hdmi_out0_driver_hdmi_phy_es0_q_m[0] + soc_hdmi_out0_driver_hdmi_phy_es0_q_m[1]) + soc_hdmi_out0_driver_hdmi_phy_es0_q_m[2]) + soc_hdmi_out0_driver_hdmi_phy_es0_q_m[3]) + soc_hdmi_out0_driver_hdmi_phy_es0_q_m[4]) + soc_hdmi_out0_driver_hdmi_phy_es0_q_m[5]) + soc_hdmi_out0_driver_hdmi_phy_es0_q_m[6]) + soc_hdmi_out0_driver_hdmi_phy_es0_q_m[7]);
	soc_hdmi_out0_driver_hdmi_phy_es0_q_m_r <= soc_hdmi_out0_driver_hdmi_phy_es0_q_m;
	soc_hdmi_out0_driver_hdmi_phy_es0_new_c0 <= soc_hdmi_out0_driver_hdmi_phy_es0_c;
	soc_hdmi_out0_driver_hdmi_phy_es0_new_de0 <= soc_hdmi_out0_driver_hdmi_phy_es0_de;
	soc_hdmi_out0_driver_hdmi_phy_es0_new_c1 <= soc_hdmi_out0_driver_hdmi_phy_es0_new_c0;
	soc_hdmi_out0_driver_hdmi_phy_es0_new_de1 <= soc_hdmi_out0_driver_hdmi_phy_es0_new_de0;
	soc_hdmi_out0_driver_hdmi_phy_es0_new_c2 <= soc_hdmi_out0_driver_hdmi_phy_es0_new_c1;
	soc_hdmi_out0_driver_hdmi_phy_es0_new_de2 <= soc_hdmi_out0_driver_hdmi_phy_es0_new_de1;
	if (soc_hdmi_out0_driver_hdmi_phy_es0_new_de2) begin
		if (((soc_hdmi_out0_driver_hdmi_phy_es0_cnt == $signed({1'd0, 1'd0})) | $signed({1'd0, (soc_hdmi_out0_driver_hdmi_phy_es0_n1q_m == soc_hdmi_out0_driver_hdmi_phy_es0_n0q_m)}))) begin
			soc_hdmi_out0_driver_hdmi_phy_es0_out[9] <= (~soc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[8]);
			soc_hdmi_out0_driver_hdmi_phy_es0_out[8] <= soc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[8];
			if (soc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[8]) begin
				soc_hdmi_out0_driver_hdmi_phy_es0_out[7:0] <= soc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[7:0];
				soc_hdmi_out0_driver_hdmi_phy_es0_cnt <= ((soc_hdmi_out0_driver_hdmi_phy_es0_cnt + $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es0_n1q_m})) - $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es0_n0q_m}));
			end else begin
				soc_hdmi_out0_driver_hdmi_phy_es0_out[7:0] <= (~soc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[7:0]);
				soc_hdmi_out0_driver_hdmi_phy_es0_cnt <= ((soc_hdmi_out0_driver_hdmi_phy_es0_cnt + $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es0_n0q_m})) - $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es0_n1q_m}));
			end
		end else begin
			if ((((~soc_hdmi_out0_driver_hdmi_phy_es0_cnt[5]) & $signed({1'd0, (soc_hdmi_out0_driver_hdmi_phy_es0_n1q_m > soc_hdmi_out0_driver_hdmi_phy_es0_n0q_m)})) | (soc_hdmi_out0_driver_hdmi_phy_es0_cnt[5] & $signed({1'd0, (soc_hdmi_out0_driver_hdmi_phy_es0_n0q_m > soc_hdmi_out0_driver_hdmi_phy_es0_n1q_m)})))) begin
				soc_hdmi_out0_driver_hdmi_phy_es0_out[9] <= 1'd1;
				soc_hdmi_out0_driver_hdmi_phy_es0_out[8] <= soc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[8];
				soc_hdmi_out0_driver_hdmi_phy_es0_out[7:0] <= (~soc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[7:0]);
				soc_hdmi_out0_driver_hdmi_phy_es0_cnt <= (((soc_hdmi_out0_driver_hdmi_phy_es0_cnt + $signed({1'd0, {soc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[8], 1'd0}})) + $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es0_n0q_m})) - $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es0_n1q_m}));
			end else begin
				soc_hdmi_out0_driver_hdmi_phy_es0_out[9] <= 1'd0;
				soc_hdmi_out0_driver_hdmi_phy_es0_out[8] <= soc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[8];
				soc_hdmi_out0_driver_hdmi_phy_es0_out[7:0] <= soc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[7:0];
				soc_hdmi_out0_driver_hdmi_phy_es0_cnt <= (((soc_hdmi_out0_driver_hdmi_phy_es0_cnt - $signed({1'd0, {(~soc_hdmi_out0_driver_hdmi_phy_es0_q_m_r[8]), 1'd0}})) + $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es0_n1q_m})) - $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es0_n0q_m}));
			end
		end
	end else begin
		soc_hdmi_out0_driver_hdmi_phy_es0_out <= vns_sync_f_array_muxed0;
		soc_hdmi_out0_driver_hdmi_phy_es0_cnt <= 1'd0;
	end
	soc_hdmi_out0_driver_hdmi_phy_es1_ce <= (~hdmi_out0_pix_rst);
	soc_hdmi_out0_driver_hdmi_phy_es1_n1d <= (((((((soc_hdmi_out0_driver_hdmi_phy_es1_d0[0] + soc_hdmi_out0_driver_hdmi_phy_es1_d0[1]) + soc_hdmi_out0_driver_hdmi_phy_es1_d0[2]) + soc_hdmi_out0_driver_hdmi_phy_es1_d0[3]) + soc_hdmi_out0_driver_hdmi_phy_es1_d0[4]) + soc_hdmi_out0_driver_hdmi_phy_es1_d0[5]) + soc_hdmi_out0_driver_hdmi_phy_es1_d0[6]) + soc_hdmi_out0_driver_hdmi_phy_es1_d0[7]);
	soc_hdmi_out0_driver_hdmi_phy_es1_d1 <= soc_hdmi_out0_driver_hdmi_phy_es1_d0;
	soc_hdmi_out0_driver_hdmi_phy_es1_q_m[0] <= soc_hdmi_out0_driver_hdmi_phy_es1_d1[0];
	soc_hdmi_out0_driver_hdmi_phy_es1_q_m[1] <= ((soc_hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es1_q_m[2] <= ((((soc_hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es1_q_m[3] <= ((((((soc_hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[3]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es1_q_m[4] <= ((((((((soc_hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[3]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[4]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es1_q_m[5] <= ((((((((((soc_hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[3]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[4]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[5]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es1_q_m[6] <= ((((((((((((soc_hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[3]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[4]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[5]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[6]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es1_q_m[7] <= ((((((((((((((soc_hdmi_out0_driver_hdmi_phy_es1_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[3]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[4]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[5]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[6]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es1_d1[7]) ^ soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es1_q_m[8] <= (~soc_hdmi_out0_driver_hdmi_phy_es1_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es1_n0q_m <= ((((((((~soc_hdmi_out0_driver_hdmi_phy_es1_q_m[0]) + (~soc_hdmi_out0_driver_hdmi_phy_es1_q_m[1])) + (~soc_hdmi_out0_driver_hdmi_phy_es1_q_m[2])) + (~soc_hdmi_out0_driver_hdmi_phy_es1_q_m[3])) + (~soc_hdmi_out0_driver_hdmi_phy_es1_q_m[4])) + (~soc_hdmi_out0_driver_hdmi_phy_es1_q_m[5])) + (~soc_hdmi_out0_driver_hdmi_phy_es1_q_m[6])) + (~soc_hdmi_out0_driver_hdmi_phy_es1_q_m[7]));
	soc_hdmi_out0_driver_hdmi_phy_es1_n1q_m <= (((((((soc_hdmi_out0_driver_hdmi_phy_es1_q_m[0] + soc_hdmi_out0_driver_hdmi_phy_es1_q_m[1]) + soc_hdmi_out0_driver_hdmi_phy_es1_q_m[2]) + soc_hdmi_out0_driver_hdmi_phy_es1_q_m[3]) + soc_hdmi_out0_driver_hdmi_phy_es1_q_m[4]) + soc_hdmi_out0_driver_hdmi_phy_es1_q_m[5]) + soc_hdmi_out0_driver_hdmi_phy_es1_q_m[6]) + soc_hdmi_out0_driver_hdmi_phy_es1_q_m[7]);
	soc_hdmi_out0_driver_hdmi_phy_es1_q_m_r <= soc_hdmi_out0_driver_hdmi_phy_es1_q_m;
	soc_hdmi_out0_driver_hdmi_phy_es1_new_c0 <= soc_hdmi_out0_driver_hdmi_phy_es1_c;
	soc_hdmi_out0_driver_hdmi_phy_es1_new_de0 <= soc_hdmi_out0_driver_hdmi_phy_es1_de;
	soc_hdmi_out0_driver_hdmi_phy_es1_new_c1 <= soc_hdmi_out0_driver_hdmi_phy_es1_new_c0;
	soc_hdmi_out0_driver_hdmi_phy_es1_new_de1 <= soc_hdmi_out0_driver_hdmi_phy_es1_new_de0;
	soc_hdmi_out0_driver_hdmi_phy_es1_new_c2 <= soc_hdmi_out0_driver_hdmi_phy_es1_new_c1;
	soc_hdmi_out0_driver_hdmi_phy_es1_new_de2 <= soc_hdmi_out0_driver_hdmi_phy_es1_new_de1;
	if (soc_hdmi_out0_driver_hdmi_phy_es1_new_de2) begin
		if (((soc_hdmi_out0_driver_hdmi_phy_es1_cnt == $signed({1'd0, 1'd0})) | $signed({1'd0, (soc_hdmi_out0_driver_hdmi_phy_es1_n1q_m == soc_hdmi_out0_driver_hdmi_phy_es1_n0q_m)}))) begin
			soc_hdmi_out0_driver_hdmi_phy_es1_out[9] <= (~soc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[8]);
			soc_hdmi_out0_driver_hdmi_phy_es1_out[8] <= soc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[8];
			if (soc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[8]) begin
				soc_hdmi_out0_driver_hdmi_phy_es1_out[7:0] <= soc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[7:0];
				soc_hdmi_out0_driver_hdmi_phy_es1_cnt <= ((soc_hdmi_out0_driver_hdmi_phy_es1_cnt + $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es1_n1q_m})) - $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es1_n0q_m}));
			end else begin
				soc_hdmi_out0_driver_hdmi_phy_es1_out[7:0] <= (~soc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[7:0]);
				soc_hdmi_out0_driver_hdmi_phy_es1_cnt <= ((soc_hdmi_out0_driver_hdmi_phy_es1_cnt + $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es1_n0q_m})) - $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es1_n1q_m}));
			end
		end else begin
			if ((((~soc_hdmi_out0_driver_hdmi_phy_es1_cnt[5]) & $signed({1'd0, (soc_hdmi_out0_driver_hdmi_phy_es1_n1q_m > soc_hdmi_out0_driver_hdmi_phy_es1_n0q_m)})) | (soc_hdmi_out0_driver_hdmi_phy_es1_cnt[5] & $signed({1'd0, (soc_hdmi_out0_driver_hdmi_phy_es1_n0q_m > soc_hdmi_out0_driver_hdmi_phy_es1_n1q_m)})))) begin
				soc_hdmi_out0_driver_hdmi_phy_es1_out[9] <= 1'd1;
				soc_hdmi_out0_driver_hdmi_phy_es1_out[8] <= soc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[8];
				soc_hdmi_out0_driver_hdmi_phy_es1_out[7:0] <= (~soc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[7:0]);
				soc_hdmi_out0_driver_hdmi_phy_es1_cnt <= (((soc_hdmi_out0_driver_hdmi_phy_es1_cnt + $signed({1'd0, {soc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[8], 1'd0}})) + $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es1_n0q_m})) - $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es1_n1q_m}));
			end else begin
				soc_hdmi_out0_driver_hdmi_phy_es1_out[9] <= 1'd0;
				soc_hdmi_out0_driver_hdmi_phy_es1_out[8] <= soc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[8];
				soc_hdmi_out0_driver_hdmi_phy_es1_out[7:0] <= soc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[7:0];
				soc_hdmi_out0_driver_hdmi_phy_es1_cnt <= (((soc_hdmi_out0_driver_hdmi_phy_es1_cnt - $signed({1'd0, {(~soc_hdmi_out0_driver_hdmi_phy_es1_q_m_r[8]), 1'd0}})) + $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es1_n1q_m})) - $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es1_n0q_m}));
			end
		end
	end else begin
		soc_hdmi_out0_driver_hdmi_phy_es1_out <= vns_sync_f_array_muxed1;
		soc_hdmi_out0_driver_hdmi_phy_es1_cnt <= 1'd0;
	end
	soc_hdmi_out0_driver_hdmi_phy_es2_ce <= (~hdmi_out0_pix_rst);
	soc_hdmi_out0_driver_hdmi_phy_es2_n1d <= (((((((soc_hdmi_out0_driver_hdmi_phy_es2_d0[0] + soc_hdmi_out0_driver_hdmi_phy_es2_d0[1]) + soc_hdmi_out0_driver_hdmi_phy_es2_d0[2]) + soc_hdmi_out0_driver_hdmi_phy_es2_d0[3]) + soc_hdmi_out0_driver_hdmi_phy_es2_d0[4]) + soc_hdmi_out0_driver_hdmi_phy_es2_d0[5]) + soc_hdmi_out0_driver_hdmi_phy_es2_d0[6]) + soc_hdmi_out0_driver_hdmi_phy_es2_d0[7]);
	soc_hdmi_out0_driver_hdmi_phy_es2_d1 <= soc_hdmi_out0_driver_hdmi_phy_es2_d0;
	soc_hdmi_out0_driver_hdmi_phy_es2_q_m[0] <= soc_hdmi_out0_driver_hdmi_phy_es2_d1[0];
	soc_hdmi_out0_driver_hdmi_phy_es2_q_m[1] <= ((soc_hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es2_q_m[2] <= ((((soc_hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es2_q_m[3] <= ((((((soc_hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[3]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es2_q_m[4] <= ((((((((soc_hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[3]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[4]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es2_q_m[5] <= ((((((((((soc_hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[3]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[4]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[5]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es2_q_m[6] <= ((((((((((((soc_hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[3]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[4]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[5]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[6]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es2_q_m[7] <= ((((((((((((((soc_hdmi_out0_driver_hdmi_phy_es2_d1[0] ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[1]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[2]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[3]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[4]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[5]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[6]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n) ^ soc_hdmi_out0_driver_hdmi_phy_es2_d1[7]) ^ soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es2_q_m[8] <= (~soc_hdmi_out0_driver_hdmi_phy_es2_q_m8_n);
	soc_hdmi_out0_driver_hdmi_phy_es2_n0q_m <= ((((((((~soc_hdmi_out0_driver_hdmi_phy_es2_q_m[0]) + (~soc_hdmi_out0_driver_hdmi_phy_es2_q_m[1])) + (~soc_hdmi_out0_driver_hdmi_phy_es2_q_m[2])) + (~soc_hdmi_out0_driver_hdmi_phy_es2_q_m[3])) + (~soc_hdmi_out0_driver_hdmi_phy_es2_q_m[4])) + (~soc_hdmi_out0_driver_hdmi_phy_es2_q_m[5])) + (~soc_hdmi_out0_driver_hdmi_phy_es2_q_m[6])) + (~soc_hdmi_out0_driver_hdmi_phy_es2_q_m[7]));
	soc_hdmi_out0_driver_hdmi_phy_es2_n1q_m <= (((((((soc_hdmi_out0_driver_hdmi_phy_es2_q_m[0] + soc_hdmi_out0_driver_hdmi_phy_es2_q_m[1]) + soc_hdmi_out0_driver_hdmi_phy_es2_q_m[2]) + soc_hdmi_out0_driver_hdmi_phy_es2_q_m[3]) + soc_hdmi_out0_driver_hdmi_phy_es2_q_m[4]) + soc_hdmi_out0_driver_hdmi_phy_es2_q_m[5]) + soc_hdmi_out0_driver_hdmi_phy_es2_q_m[6]) + soc_hdmi_out0_driver_hdmi_phy_es2_q_m[7]);
	soc_hdmi_out0_driver_hdmi_phy_es2_q_m_r <= soc_hdmi_out0_driver_hdmi_phy_es2_q_m;
	soc_hdmi_out0_driver_hdmi_phy_es2_new_c0 <= soc_hdmi_out0_driver_hdmi_phy_es2_c;
	soc_hdmi_out0_driver_hdmi_phy_es2_new_de0 <= soc_hdmi_out0_driver_hdmi_phy_es2_de;
	soc_hdmi_out0_driver_hdmi_phy_es2_new_c1 <= soc_hdmi_out0_driver_hdmi_phy_es2_new_c0;
	soc_hdmi_out0_driver_hdmi_phy_es2_new_de1 <= soc_hdmi_out0_driver_hdmi_phy_es2_new_de0;
	soc_hdmi_out0_driver_hdmi_phy_es2_new_c2 <= soc_hdmi_out0_driver_hdmi_phy_es2_new_c1;
	soc_hdmi_out0_driver_hdmi_phy_es2_new_de2 <= soc_hdmi_out0_driver_hdmi_phy_es2_new_de1;
	if (soc_hdmi_out0_driver_hdmi_phy_es2_new_de2) begin
		if (((soc_hdmi_out0_driver_hdmi_phy_es2_cnt == $signed({1'd0, 1'd0})) | $signed({1'd0, (soc_hdmi_out0_driver_hdmi_phy_es2_n1q_m == soc_hdmi_out0_driver_hdmi_phy_es2_n0q_m)}))) begin
			soc_hdmi_out0_driver_hdmi_phy_es2_out[9] <= (~soc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[8]);
			soc_hdmi_out0_driver_hdmi_phy_es2_out[8] <= soc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[8];
			if (soc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[8]) begin
				soc_hdmi_out0_driver_hdmi_phy_es2_out[7:0] <= soc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[7:0];
				soc_hdmi_out0_driver_hdmi_phy_es2_cnt <= ((soc_hdmi_out0_driver_hdmi_phy_es2_cnt + $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es2_n1q_m})) - $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es2_n0q_m}));
			end else begin
				soc_hdmi_out0_driver_hdmi_phy_es2_out[7:0] <= (~soc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[7:0]);
				soc_hdmi_out0_driver_hdmi_phy_es2_cnt <= ((soc_hdmi_out0_driver_hdmi_phy_es2_cnt + $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es2_n0q_m})) - $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es2_n1q_m}));
			end
		end else begin
			if ((((~soc_hdmi_out0_driver_hdmi_phy_es2_cnt[5]) & $signed({1'd0, (soc_hdmi_out0_driver_hdmi_phy_es2_n1q_m > soc_hdmi_out0_driver_hdmi_phy_es2_n0q_m)})) | (soc_hdmi_out0_driver_hdmi_phy_es2_cnt[5] & $signed({1'd0, (soc_hdmi_out0_driver_hdmi_phy_es2_n0q_m > soc_hdmi_out0_driver_hdmi_phy_es2_n1q_m)})))) begin
				soc_hdmi_out0_driver_hdmi_phy_es2_out[9] <= 1'd1;
				soc_hdmi_out0_driver_hdmi_phy_es2_out[8] <= soc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[8];
				soc_hdmi_out0_driver_hdmi_phy_es2_out[7:0] <= (~soc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[7:0]);
				soc_hdmi_out0_driver_hdmi_phy_es2_cnt <= (((soc_hdmi_out0_driver_hdmi_phy_es2_cnt + $signed({1'd0, {soc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[8], 1'd0}})) + $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es2_n0q_m})) - $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es2_n1q_m}));
			end else begin
				soc_hdmi_out0_driver_hdmi_phy_es2_out[9] <= 1'd0;
				soc_hdmi_out0_driver_hdmi_phy_es2_out[8] <= soc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[8];
				soc_hdmi_out0_driver_hdmi_phy_es2_out[7:0] <= soc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[7:0];
				soc_hdmi_out0_driver_hdmi_phy_es2_cnt <= (((soc_hdmi_out0_driver_hdmi_phy_es2_cnt - $signed({1'd0, {(~soc_hdmi_out0_driver_hdmi_phy_es2_q_m_r[8]), 1'd0}})) + $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es2_n1q_m})) - $signed({1'd0, soc_hdmi_out0_driver_hdmi_phy_es2_n0q_m}));
			end
		end
	end else begin
		soc_hdmi_out0_driver_hdmi_phy_es2_out <= vns_sync_f_array_muxed2;
		soc_hdmi_out0_driver_hdmi_phy_es2_cnt <= 1'd0;
	end
	if (hdmi_out0_pix_rst) begin
		soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q <= 3'd0;
		soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q_binary <= 3'd0;
		soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q <= 5'd0;
		soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q_binary <= 5'd0;
		soc_hdmi_out0_dram_port_cmd_buffer_level <= 3'd0;
		soc_hdmi_out0_dram_port_cmd_buffer_produce <= 2'd0;
		soc_hdmi_out0_dram_port_cmd_buffer_consume <= 2'd0;
		soc_hdmi_out0_dram_port_counter <= 3'd0;
		soc_hdmi_out0_dram_port_rdata_buffer_valid_n <= 1'd0;
		soc_hdmi_out0_dram_port_rdata_buffer_first_n <= 1'd0;
		soc_hdmi_out0_dram_port_rdata_buffer_last_n <= 1'd0;
		soc_hdmi_out0_dram_port_rdata_converter_converter_mux <= 3'd0;
		soc_hdmi_out0_dram_port_rdata_chunk <= 8'd1;
		soc_hdmi_out0_core_underflow_counter_status <= 32'd0;
		soc_hdmi_out0_core_initiator_cdc_graycounter1_q <= 2'd0;
		soc_hdmi_out0_core_initiator_cdc_graycounter1_q_binary <= 2'd0;
		soc_hdmi_out0_core_timinggenerator_source_last <= 1'd0;
		soc_hdmi_out0_core_timinggenerator_hactive <= 1'd0;
		soc_hdmi_out0_core_timinggenerator_vactive <= 1'd0;
		soc_hdmi_out0_core_timinggenerator_hcounter <= 12'd0;
		soc_hdmi_out0_core_timinggenerator_vcounter <= 12'd0;
		soc_hdmi_out0_core_dmareader_rsv_level <= 13'd0;
		soc_hdmi_out0_core_dmareader_fifo_readable <= 1'd0;
		soc_hdmi_out0_core_dmareader_fifo_level0 <= 13'd0;
		soc_hdmi_out0_core_dmareader_fifo_produce <= 12'd0;
		soc_hdmi_out0_core_dmareader_fifo_consume <= 12'd0;
		soc_hdmi_out0_core_dmareader_offset <= 28'd0;
		soc_hdmi_out0_core_underflow_counter <= 32'd0;
		soc_hdmi_out0_driver_s7hdmioutclocking_ce <= 1'd0;
		soc_hdmi_out0_driver_hdmi_phy_es0_out <= 10'd0;
		soc_hdmi_out0_driver_hdmi_phy_es0_d1 <= 8'd0;
		soc_hdmi_out0_driver_hdmi_phy_es0_n1d <= 4'd0;
		soc_hdmi_out0_driver_hdmi_phy_es0_q_m <= 9'd0;
		soc_hdmi_out0_driver_hdmi_phy_es0_q_m_r <= 9'd0;
		soc_hdmi_out0_driver_hdmi_phy_es0_n0q_m <= 4'd0;
		soc_hdmi_out0_driver_hdmi_phy_es0_n1q_m <= 4'd0;
		soc_hdmi_out0_driver_hdmi_phy_es0_cnt <= 6'sd64;
		soc_hdmi_out0_driver_hdmi_phy_es0_new_c0 <= 2'd0;
		soc_hdmi_out0_driver_hdmi_phy_es0_new_de0 <= 1'd0;
		soc_hdmi_out0_driver_hdmi_phy_es0_new_c1 <= 2'd0;
		soc_hdmi_out0_driver_hdmi_phy_es0_new_de1 <= 1'd0;
		soc_hdmi_out0_driver_hdmi_phy_es0_new_c2 <= 2'd0;
		soc_hdmi_out0_driver_hdmi_phy_es0_new_de2 <= 1'd0;
		soc_hdmi_out0_driver_hdmi_phy_es0_ce <= 1'd0;
		soc_hdmi_out0_driver_hdmi_phy_es1_out <= 10'd0;
		soc_hdmi_out0_driver_hdmi_phy_es1_d1 <= 8'd0;
		soc_hdmi_out0_driver_hdmi_phy_es1_n1d <= 4'd0;
		soc_hdmi_out0_driver_hdmi_phy_es1_q_m <= 9'd0;
		soc_hdmi_out0_driver_hdmi_phy_es1_q_m_r <= 9'd0;
		soc_hdmi_out0_driver_hdmi_phy_es1_n0q_m <= 4'd0;
		soc_hdmi_out0_driver_hdmi_phy_es1_n1q_m <= 4'd0;
		soc_hdmi_out0_driver_hdmi_phy_es1_cnt <= 6'sd64;
		soc_hdmi_out0_driver_hdmi_phy_es1_new_c0 <= 2'd0;
		soc_hdmi_out0_driver_hdmi_phy_es1_new_de0 <= 1'd0;
		soc_hdmi_out0_driver_hdmi_phy_es1_new_c1 <= 2'd0;
		soc_hdmi_out0_driver_hdmi_phy_es1_new_de1 <= 1'd0;
		soc_hdmi_out0_driver_hdmi_phy_es1_new_c2 <= 2'd0;
		soc_hdmi_out0_driver_hdmi_phy_es1_new_de2 <= 1'd0;
		soc_hdmi_out0_driver_hdmi_phy_es1_ce <= 1'd0;
		soc_hdmi_out0_driver_hdmi_phy_es2_out <= 10'd0;
		soc_hdmi_out0_driver_hdmi_phy_es2_d1 <= 8'd0;
		soc_hdmi_out0_driver_hdmi_phy_es2_n1d <= 4'd0;
		soc_hdmi_out0_driver_hdmi_phy_es2_q_m <= 9'd0;
		soc_hdmi_out0_driver_hdmi_phy_es2_q_m_r <= 9'd0;
		soc_hdmi_out0_driver_hdmi_phy_es2_n0q_m <= 4'd0;
		soc_hdmi_out0_driver_hdmi_phy_es2_n1q_m <= 4'd0;
		soc_hdmi_out0_driver_hdmi_phy_es2_cnt <= 6'sd64;
		soc_hdmi_out0_driver_hdmi_phy_es2_new_c0 <= 2'd0;
		soc_hdmi_out0_driver_hdmi_phy_es2_new_de0 <= 1'd0;
		soc_hdmi_out0_driver_hdmi_phy_es2_new_c1 <= 2'd0;
		soc_hdmi_out0_driver_hdmi_phy_es2_new_de1 <= 1'd0;
		soc_hdmi_out0_driver_hdmi_phy_es2_new_c2 <= 2'd0;
		soc_hdmi_out0_driver_hdmi_phy_es2_new_de2 <= 1'd0;
		soc_hdmi_out0_driver_hdmi_phy_es2_ce <= 1'd0;
		soc_hdmi_out0_resetinserter_y_fifo_level <= 3'd0;
		soc_hdmi_out0_resetinserter_y_fifo_produce <= 2'd0;
		soc_hdmi_out0_resetinserter_y_fifo_consume <= 2'd0;
		soc_hdmi_out0_resetinserter_cb_fifo_level <= 3'd0;
		soc_hdmi_out0_resetinserter_cb_fifo_produce <= 2'd0;
		soc_hdmi_out0_resetinserter_cb_fifo_consume <= 2'd0;
		soc_hdmi_out0_resetinserter_cr_fifo_level <= 3'd0;
		soc_hdmi_out0_resetinserter_cr_fifo_produce <= 2'd0;
		soc_hdmi_out0_resetinserter_cr_fifo_consume <= 2'd0;
		soc_hdmi_out0_resetinserter_parity_in <= 1'd0;
		soc_hdmi_out0_resetinserter_parity_out <= 1'd0;
		soc_hdmi_out0_source_r <= 8'd0;
		soc_hdmi_out0_source_g <= 8'd0;
		soc_hdmi_out0_source_b <= 8'd0;
		soc_hdmi_out0_record0_ycbcr_n_y <= 8'd0;
		soc_hdmi_out0_record0_ycbcr_n_cb <= 8'd0;
		soc_hdmi_out0_record0_ycbcr_n_cr <= 8'd0;
		soc_hdmi_out0_record1_ycbcr_n_y <= 8'd0;
		soc_hdmi_out0_record1_ycbcr_n_cb <= 8'd0;
		soc_hdmi_out0_record1_ycbcr_n_cr <= 8'd0;
		soc_hdmi_out0_record2_ycbcr_n_y <= 8'd0;
		soc_hdmi_out0_record2_ycbcr_n_cb <= 8'd0;
		soc_hdmi_out0_record2_ycbcr_n_cr <= 8'd0;
		soc_hdmi_out0_record3_ycbcr_n_y <= 8'd0;
		soc_hdmi_out0_record3_ycbcr_n_cb <= 8'd0;
		soc_hdmi_out0_record3_ycbcr_n_cr <= 8'd0;
		soc_hdmi_out0_cb_minus_coffset <= 9'sd512;
		soc_hdmi_out0_cr_minus_coffset <= 9'sd512;
		soc_hdmi_out0_y_minus_yoffset <= 9'sd512;
		soc_hdmi_out0_cr_minus_coffset_mult_acoef <= 20'sd1048576;
		soc_hdmi_out0_cb_minus_coffset_mult_bcoef <= 20'sd1048576;
		soc_hdmi_out0_cr_minus_coffset_mult_ccoef <= 20'sd1048576;
		soc_hdmi_out0_cb_minus_coffset_mult_dcoef <= 20'sd1048576;
		soc_hdmi_out0_r <= 12'sd4096;
		soc_hdmi_out0_g <= 12'sd4096;
		soc_hdmi_out0_b <= 12'sd4096;
		soc_hdmi_out0_valid_n0 <= 1'd0;
		soc_hdmi_out0_valid_n1 <= 1'd0;
		soc_hdmi_out0_valid_n2 <= 1'd0;
		soc_hdmi_out0_valid_n3 <= 1'd0;
		soc_hdmi_out0_first_n0 <= 1'd0;
		soc_hdmi_out0_last_n0 <= 1'd0;
		soc_hdmi_out0_first_n1 <= 1'd0;
		soc_hdmi_out0_last_n1 <= 1'd0;
		soc_hdmi_out0_first_n2 <= 1'd0;
		soc_hdmi_out0_last_n2 <= 1'd0;
		soc_hdmi_out0_first_n3 <= 1'd0;
		soc_hdmi_out0_last_n3 <= 1'd0;
		soc_hdmi_out0_next_s0 <= 1'd0;
		soc_hdmi_out0_next_s1 <= 1'd0;
		soc_hdmi_out0_next_s2 <= 1'd0;
		soc_hdmi_out0_next_s3 <= 1'd0;
		soc_hdmi_out0_next_s4 <= 1'd0;
		soc_hdmi_out0_next_s5 <= 1'd0;
		soc_hdmi_out0_next_s6 <= 1'd0;
		soc_hdmi_out0_next_s7 <= 1'd0;
		soc_hdmi_out0_next_s8 <= 1'd0;
		soc_hdmi_out0_next_s9 <= 1'd0;
		soc_hdmi_out0_next_s10 <= 1'd0;
		soc_hdmi_out0_next_s11 <= 1'd0;
		soc_hdmi_out0_next_s12 <= 1'd0;
		soc_hdmi_out0_next_s13 <= 1'd0;
		soc_hdmi_out0_next_s14 <= 1'd0;
		soc_hdmi_out0_next_s15 <= 1'd0;
		soc_hdmi_out0_next_s16 <= 1'd0;
		soc_hdmi_out0_next_s17 <= 1'd0;
		soc_hdmi_out0_de_r <= 1'd0;
		soc_hdmi_out0_core_source_valid_d <= 1'd0;
		soc_hdmi_out0_core_source_data_d <= 16'd0;
		vns_videoout_state <= 1'd0;
	end
	vns_xilinxmultiregimpl49_regs0 <= soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q;
	vns_xilinxmultiregimpl49_regs1 <= vns_xilinxmultiregimpl49_regs0;
	vns_xilinxmultiregimpl50_regs0 <= soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q;
	vns_xilinxmultiregimpl50_regs1 <= vns_xilinxmultiregimpl50_regs0;
	vns_xilinxmultiregimpl52_regs0 <= soc_hdmi_out0_core_initiator_cdc_graycounter0_q;
	vns_xilinxmultiregimpl52_regs1 <= vns_xilinxmultiregimpl52_regs0;
	vns_xilinxmultiregimpl55_regs0 <= soc_hdmi_out0_core_toggle_i;
	vns_xilinxmultiregimpl55_regs1 <= vns_xilinxmultiregimpl55_regs0;
end

always @(posedge pix1p25x_clk) begin
	if (soc_s7datacapture0_reset_lateness) begin
		soc_s7datacapture0_lateness <= 8'd128;
	end else begin
		if (((~soc_s7datacapture0_too_late) & (~soc_s7datacapture0_too_early))) begin
			if (soc_s7datacapture0_dec) begin
				soc_s7datacapture0_lateness <= (soc_s7datacapture0_lateness + 1'd1);
			end
			if (soc_s7datacapture0_inc) begin
				soc_s7datacapture0_lateness <= (soc_s7datacapture0_lateness - 1'd1);
			end
		end
	end
	soc_s7datacapture0_mdata_d <= soc_s7datacapture0_mdata;
	soc_s7datacapture0_do_delay_rst_toggle_o_r <= soc_s7datacapture0_do_delay_rst_toggle_o;
	soc_s7datacapture0_do_delay_master_inc_toggle_o_r <= soc_s7datacapture0_do_delay_master_inc_toggle_o;
	soc_s7datacapture0_do_delay_master_dec_toggle_o_r <= soc_s7datacapture0_do_delay_master_dec_toggle_o;
	soc_s7datacapture0_do_delay_slave_inc_toggle_o_r <= soc_s7datacapture0_do_delay_slave_inc_toggle_o;
	soc_s7datacapture0_do_delay_slave_dec_toggle_o_r <= soc_s7datacapture0_do_delay_slave_dec_toggle_o;
	soc_s7datacapture0_do_reset_lateness_toggle_o_r <= soc_s7datacapture0_do_reset_lateness_toggle_o;
	if (soc_s7datacapture1_reset_lateness) begin
		soc_s7datacapture1_lateness <= 8'd128;
	end else begin
		if (((~soc_s7datacapture1_too_late) & (~soc_s7datacapture1_too_early))) begin
			if (soc_s7datacapture1_dec) begin
				soc_s7datacapture1_lateness <= (soc_s7datacapture1_lateness + 1'd1);
			end
			if (soc_s7datacapture1_inc) begin
				soc_s7datacapture1_lateness <= (soc_s7datacapture1_lateness - 1'd1);
			end
		end
	end
	soc_s7datacapture1_mdata_d <= soc_s7datacapture1_mdata;
	soc_s7datacapture1_do_delay_rst_toggle_o_r <= soc_s7datacapture1_do_delay_rst_toggle_o;
	soc_s7datacapture1_do_delay_master_inc_toggle_o_r <= soc_s7datacapture1_do_delay_master_inc_toggle_o;
	soc_s7datacapture1_do_delay_master_dec_toggle_o_r <= soc_s7datacapture1_do_delay_master_dec_toggle_o;
	soc_s7datacapture1_do_delay_slave_inc_toggle_o_r <= soc_s7datacapture1_do_delay_slave_inc_toggle_o;
	soc_s7datacapture1_do_delay_slave_dec_toggle_o_r <= soc_s7datacapture1_do_delay_slave_dec_toggle_o;
	soc_s7datacapture1_do_reset_lateness_toggle_o_r <= soc_s7datacapture1_do_reset_lateness_toggle_o;
	if (soc_s7datacapture2_reset_lateness) begin
		soc_s7datacapture2_lateness <= 8'd128;
	end else begin
		if (((~soc_s7datacapture2_too_late) & (~soc_s7datacapture2_too_early))) begin
			if (soc_s7datacapture2_dec) begin
				soc_s7datacapture2_lateness <= (soc_s7datacapture2_lateness + 1'd1);
			end
			if (soc_s7datacapture2_inc) begin
				soc_s7datacapture2_lateness <= (soc_s7datacapture2_lateness - 1'd1);
			end
		end
	end
	soc_s7datacapture2_mdata_d <= soc_s7datacapture2_mdata;
	soc_s7datacapture2_do_delay_rst_toggle_o_r <= soc_s7datacapture2_do_delay_rst_toggle_o;
	soc_s7datacapture2_do_delay_master_inc_toggle_o_r <= soc_s7datacapture2_do_delay_master_inc_toggle_o;
	soc_s7datacapture2_do_delay_master_dec_toggle_o_r <= soc_s7datacapture2_do_delay_master_dec_toggle_o;
	soc_s7datacapture2_do_delay_slave_inc_toggle_o_r <= soc_s7datacapture2_do_delay_slave_inc_toggle_o;
	soc_s7datacapture2_do_delay_slave_dec_toggle_o_r <= soc_s7datacapture2_do_delay_slave_dec_toggle_o;
	soc_s7datacapture2_do_reset_lateness_toggle_o_r <= soc_s7datacapture2_do_reset_lateness_toggle_o;
	if (pix1p25x_rst) begin
		soc_s7datacapture0_mdata_d <= 8'd0;
		soc_s7datacapture0_lateness <= 8'd128;
		soc_s7datacapture1_mdata_d <= 8'd0;
		soc_s7datacapture1_lateness <= 8'd128;
		soc_s7datacapture2_mdata_d <= 8'd0;
		soc_s7datacapture2_lateness <= 8'd128;
	end
	vns_xilinxmultiregimpl9_regs0 <= soc_s7datacapture0_do_delay_rst_toggle_i;
	vns_xilinxmultiregimpl9_regs1 <= vns_xilinxmultiregimpl9_regs0;
	vns_xilinxmultiregimpl10_regs0 <= soc_s7datacapture0_do_delay_master_inc_toggle_i;
	vns_xilinxmultiregimpl10_regs1 <= vns_xilinxmultiregimpl10_regs0;
	vns_xilinxmultiregimpl11_regs0 <= soc_s7datacapture0_do_delay_master_dec_toggle_i;
	vns_xilinxmultiregimpl11_regs1 <= vns_xilinxmultiregimpl11_regs0;
	vns_xilinxmultiregimpl12_regs0 <= soc_s7datacapture0_do_delay_slave_inc_toggle_i;
	vns_xilinxmultiregimpl12_regs1 <= vns_xilinxmultiregimpl12_regs0;
	vns_xilinxmultiregimpl13_regs0 <= soc_s7datacapture0_do_delay_slave_dec_toggle_i;
	vns_xilinxmultiregimpl13_regs1 <= vns_xilinxmultiregimpl13_regs0;
	vns_xilinxmultiregimpl15_regs0 <= soc_s7datacapture0_do_reset_lateness_toggle_i;
	vns_xilinxmultiregimpl15_regs1 <= vns_xilinxmultiregimpl15_regs0;
	vns_xilinxmultiregimpl19_regs0 <= soc_s7datacapture1_do_delay_rst_toggle_i;
	vns_xilinxmultiregimpl19_regs1 <= vns_xilinxmultiregimpl19_regs0;
	vns_xilinxmultiregimpl20_regs0 <= soc_s7datacapture1_do_delay_master_inc_toggle_i;
	vns_xilinxmultiregimpl20_regs1 <= vns_xilinxmultiregimpl20_regs0;
	vns_xilinxmultiregimpl21_regs0 <= soc_s7datacapture1_do_delay_master_dec_toggle_i;
	vns_xilinxmultiregimpl21_regs1 <= vns_xilinxmultiregimpl21_regs0;
	vns_xilinxmultiregimpl22_regs0 <= soc_s7datacapture1_do_delay_slave_inc_toggle_i;
	vns_xilinxmultiregimpl22_regs1 <= vns_xilinxmultiregimpl22_regs0;
	vns_xilinxmultiregimpl23_regs0 <= soc_s7datacapture1_do_delay_slave_dec_toggle_i;
	vns_xilinxmultiregimpl23_regs1 <= vns_xilinxmultiregimpl23_regs0;
	vns_xilinxmultiregimpl25_regs0 <= soc_s7datacapture1_do_reset_lateness_toggle_i;
	vns_xilinxmultiregimpl25_regs1 <= vns_xilinxmultiregimpl25_regs0;
	vns_xilinxmultiregimpl29_regs0 <= soc_s7datacapture2_do_delay_rst_toggle_i;
	vns_xilinxmultiregimpl29_regs1 <= vns_xilinxmultiregimpl29_regs0;
	vns_xilinxmultiregimpl30_regs0 <= soc_s7datacapture2_do_delay_master_inc_toggle_i;
	vns_xilinxmultiregimpl30_regs1 <= vns_xilinxmultiregimpl30_regs0;
	vns_xilinxmultiregimpl31_regs0 <= soc_s7datacapture2_do_delay_master_dec_toggle_i;
	vns_xilinxmultiregimpl31_regs1 <= vns_xilinxmultiregimpl31_regs0;
	vns_xilinxmultiregimpl32_regs0 <= soc_s7datacapture2_do_delay_slave_inc_toggle_i;
	vns_xilinxmultiregimpl32_regs1 <= vns_xilinxmultiregimpl32_regs0;
	vns_xilinxmultiregimpl33_regs0 <= soc_s7datacapture2_do_delay_slave_dec_toggle_i;
	vns_xilinxmultiregimpl33_regs1 <= vns_xilinxmultiregimpl33_regs0;
	vns_xilinxmultiregimpl35_regs0 <= soc_s7datacapture2_do_reset_lateness_toggle_i;
	vns_xilinxmultiregimpl35_regs1 <= vns_xilinxmultiregimpl35_regs0;
end

always @(posedge sys_clk) begin
	soc_videosoc_videosoc_rom_bus_ack <= 1'd0;
	if (((soc_videosoc_videosoc_rom_bus_cyc & soc_videosoc_videosoc_rom_bus_stb) & (~soc_videosoc_videosoc_rom_bus_ack))) begin
		soc_videosoc_videosoc_rom_bus_ack <= 1'd1;
	end
	soc_videosoc_videosoc_sram_bus_ack <= 1'd0;
	if (((soc_videosoc_videosoc_sram_bus_cyc & soc_videosoc_videosoc_sram_bus_stb) & (~soc_videosoc_videosoc_sram_bus_ack))) begin
		soc_videosoc_videosoc_sram_bus_ack <= 1'd1;
	end
	soc_videosoc_videosoc_interface_we <= 1'd0;
	soc_videosoc_videosoc_interface_dat_w <= soc_videosoc_videosoc_bus_wishbone_dat_w;
	soc_videosoc_videosoc_interface_adr <= soc_videosoc_videosoc_bus_wishbone_adr;
	soc_videosoc_videosoc_bus_wishbone_dat_r <= soc_videosoc_videosoc_interface_dat_r;
	if ((soc_videosoc_videosoc_counter == 1'd1)) begin
		soc_videosoc_videosoc_interface_we <= soc_videosoc_videosoc_bus_wishbone_we;
	end
	if ((soc_videosoc_videosoc_counter == 2'd2)) begin
		soc_videosoc_videosoc_bus_wishbone_ack <= 1'd1;
	end
	if ((soc_videosoc_videosoc_counter == 2'd3)) begin
		soc_videosoc_videosoc_bus_wishbone_ack <= 1'd0;
	end
	if ((soc_videosoc_videosoc_counter != 1'd0)) begin
		soc_videosoc_videosoc_counter <= (soc_videosoc_videosoc_counter + 1'd1);
	end else begin
		if ((soc_videosoc_videosoc_bus_wishbone_cyc & soc_videosoc_videosoc_bus_wishbone_stb)) begin
			soc_videosoc_videosoc_counter <= 1'd1;
		end
	end
	if (soc_videosoc_videosoc_en_storage) begin
		if ((soc_videosoc_videosoc_value == 1'd0)) begin
			soc_videosoc_videosoc_value <= soc_videosoc_videosoc_reload_storage;
		end else begin
			soc_videosoc_videosoc_value <= (soc_videosoc_videosoc_value - 1'd1);
		end
	end else begin
		soc_videosoc_videosoc_value <= soc_videosoc_videosoc_load_storage;
	end
	if (soc_videosoc_videosoc_update_value_re) begin
		soc_videosoc_videosoc_value_status <= soc_videosoc_videosoc_value;
	end
	if (soc_videosoc_videosoc_zero_clear) begin
		soc_videosoc_videosoc_zero_pending <= 1'd0;
	end
	soc_videosoc_videosoc_zero_old_trigger <= soc_videosoc_videosoc_zero_trigger;
	if (((~soc_videosoc_videosoc_zero_trigger) & soc_videosoc_videosoc_zero_old_trigger)) begin
		soc_videosoc_videosoc_zero_pending <= 1'd1;
	end
	if (soc_videosoc_uart_tx_clear) begin
		soc_videosoc_uart_tx_pending <= 1'd0;
	end
	soc_videosoc_uart_tx_old_trigger <= soc_videosoc_uart_tx_trigger;
	if (((~soc_videosoc_uart_tx_trigger) & soc_videosoc_uart_tx_old_trigger)) begin
		soc_videosoc_uart_tx_pending <= 1'd1;
	end
	if (soc_videosoc_uart_rx_clear) begin
		soc_videosoc_uart_rx_pending <= 1'd0;
	end
	soc_videosoc_uart_rx_old_trigger <= soc_videosoc_uart_rx_trigger;
	if (((~soc_videosoc_uart_rx_trigger) & soc_videosoc_uart_rx_old_trigger)) begin
		soc_videosoc_uart_rx_pending <= 1'd1;
	end
	if (((soc_videosoc_uart_tx_fifo_syncfifo_we & soc_videosoc_uart_tx_fifo_syncfifo_writable) & (~soc_videosoc_uart_tx_fifo_replace))) begin
		soc_videosoc_uart_tx_fifo_produce <= (soc_videosoc_uart_tx_fifo_produce + 1'd1);
	end
	if (soc_videosoc_uart_tx_fifo_do_read) begin
		soc_videosoc_uart_tx_fifo_consume <= (soc_videosoc_uart_tx_fifo_consume + 1'd1);
	end
	if (((soc_videosoc_uart_tx_fifo_syncfifo_we & soc_videosoc_uart_tx_fifo_syncfifo_writable) & (~soc_videosoc_uart_tx_fifo_replace))) begin
		if ((~soc_videosoc_uart_tx_fifo_do_read)) begin
			soc_videosoc_uart_tx_fifo_level <= (soc_videosoc_uart_tx_fifo_level + 1'd1);
		end
	end else begin
		if (soc_videosoc_uart_tx_fifo_do_read) begin
			soc_videosoc_uart_tx_fifo_level <= (soc_videosoc_uart_tx_fifo_level - 1'd1);
		end
	end
	if (((soc_videosoc_uart_rx_fifo_syncfifo_we & soc_videosoc_uart_rx_fifo_syncfifo_writable) & (~soc_videosoc_uart_rx_fifo_replace))) begin
		soc_videosoc_uart_rx_fifo_produce <= (soc_videosoc_uart_rx_fifo_produce + 1'd1);
	end
	if (soc_videosoc_uart_rx_fifo_do_read) begin
		soc_videosoc_uart_rx_fifo_consume <= (soc_videosoc_uart_rx_fifo_consume + 1'd1);
	end
	if (((soc_videosoc_uart_rx_fifo_syncfifo_we & soc_videosoc_uart_rx_fifo_syncfifo_writable) & (~soc_videosoc_uart_rx_fifo_replace))) begin
		if ((~soc_videosoc_uart_rx_fifo_do_read)) begin
			soc_videosoc_uart_rx_fifo_level <= (soc_videosoc_uart_rx_fifo_level + 1'd1);
		end
	end else begin
		if (soc_videosoc_uart_rx_fifo_do_read) begin
			soc_videosoc_uart_rx_fifo_level <= (soc_videosoc_uart_rx_fifo_level - 1'd1);
		end
	end
	if (soc_videosoc_bridge_byte_counter_reset) begin
		soc_videosoc_bridge_byte_counter <= 1'd0;
	end else begin
		if (soc_videosoc_bridge_byte_counter_ce) begin
			soc_videosoc_bridge_byte_counter <= (soc_videosoc_bridge_byte_counter + 1'd1);
		end
	end
	if (soc_videosoc_bridge_word_counter_reset) begin
		soc_videosoc_bridge_word_counter <= 1'd0;
	end else begin
		if (soc_videosoc_bridge_word_counter_ce) begin
			soc_videosoc_bridge_word_counter <= (soc_videosoc_bridge_word_counter + 1'd1);
		end
	end
	if (soc_videosoc_bridge_cmd_ce) begin
		soc_videosoc_bridge_cmd <= soc_videosoc_rs232phyinterface1_source_payload_data;
	end
	if (soc_videosoc_bridge_length_ce) begin
		soc_videosoc_bridge_length <= soc_videosoc_rs232phyinterface1_source_payload_data;
	end
	if (soc_videosoc_bridge_address_ce) begin
		soc_videosoc_bridge_address <= {soc_videosoc_bridge_address[23:0], soc_videosoc_rs232phyinterface1_source_payload_data};
	end
	if (soc_videosoc_bridge_rx_data_ce) begin
		soc_videosoc_bridge_data <= {soc_videosoc_bridge_data[23:0], soc_videosoc_rs232phyinterface1_source_payload_data};
	end else begin
		if (soc_videosoc_bridge_tx_data_ce) begin
			soc_videosoc_bridge_data <= soc_videosoc_bridge_wishbone_dat_r;
		end
	end
	vns_wishbonestreamingbridge_state <= vns_wishbonestreamingbridge_next_state;
	if (soc_videosoc_bridge_reset) begin
		vns_wishbonestreamingbridge_state <= 3'd0;
	end
	if (soc_videosoc_bridge_wait) begin
		if ((~soc_videosoc_bridge_done)) begin
			soc_videosoc_bridge_count <= (soc_videosoc_bridge_count - 1'd1);
		end
	end else begin
		soc_videosoc_bridge_count <= 24'd10000000;
	end
	soc_videosoc_uart_phy_sink_ready <= 1'd0;
	if (((soc_videosoc_uart_phy_sink_valid & (~soc_videosoc_uart_phy_tx_busy)) & (~soc_videosoc_uart_phy_sink_ready))) begin
		soc_videosoc_uart_phy_tx_reg <= soc_videosoc_uart_phy_sink_payload_data;
		soc_videosoc_uart_phy_tx_bitcount <= 1'd0;
		soc_videosoc_uart_phy_tx_busy <= 1'd1;
		serial_tx <= 1'd0;
	end else begin
		if ((soc_videosoc_uart_phy_uart_clk_txen & soc_videosoc_uart_phy_tx_busy)) begin
			soc_videosoc_uart_phy_tx_bitcount <= (soc_videosoc_uart_phy_tx_bitcount + 1'd1);
			if ((soc_videosoc_uart_phy_tx_bitcount == 4'd8)) begin
				serial_tx <= 1'd1;
			end else begin
				if ((soc_videosoc_uart_phy_tx_bitcount == 4'd9)) begin
					serial_tx <= 1'd1;
					soc_videosoc_uart_phy_tx_busy <= 1'd0;
					soc_videosoc_uart_phy_sink_ready <= 1'd1;
				end else begin
					serial_tx <= soc_videosoc_uart_phy_tx_reg[0];
					soc_videosoc_uart_phy_tx_reg <= {1'd0, soc_videosoc_uart_phy_tx_reg[7:1]};
				end
			end
		end
	end
	if (soc_videosoc_uart_phy_tx_busy) begin
		{soc_videosoc_uart_phy_uart_clk_txen, soc_videosoc_uart_phy_phase_accumulator_tx} <= (soc_videosoc_uart_phy_phase_accumulator_tx + soc_videosoc_uart_phy_storage);
	end else begin
		{soc_videosoc_uart_phy_uart_clk_txen, soc_videosoc_uart_phy_phase_accumulator_tx} <= 1'd0;
	end
	soc_videosoc_uart_phy_source_valid <= 1'd0;
	soc_videosoc_uart_phy_rx_r <= soc_videosoc_uart_phy_rx;
	if ((~soc_videosoc_uart_phy_rx_busy)) begin
		if (((~soc_videosoc_uart_phy_rx) & soc_videosoc_uart_phy_rx_r)) begin
			soc_videosoc_uart_phy_rx_busy <= 1'd1;
			soc_videosoc_uart_phy_rx_bitcount <= 1'd0;
		end
	end else begin
		if (soc_videosoc_uart_phy_uart_clk_rxen) begin
			soc_videosoc_uart_phy_rx_bitcount <= (soc_videosoc_uart_phy_rx_bitcount + 1'd1);
			if ((soc_videosoc_uart_phy_rx_bitcount == 1'd0)) begin
				if (soc_videosoc_uart_phy_rx) begin
					soc_videosoc_uart_phy_rx_busy <= 1'd0;
				end
			end else begin
				if ((soc_videosoc_uart_phy_rx_bitcount == 4'd9)) begin
					soc_videosoc_uart_phy_rx_busy <= 1'd0;
					if (soc_videosoc_uart_phy_rx) begin
						soc_videosoc_uart_phy_source_payload_data <= soc_videosoc_uart_phy_rx_reg;
						soc_videosoc_uart_phy_source_valid <= 1'd1;
					end
				end else begin
					soc_videosoc_uart_phy_rx_reg <= {soc_videosoc_uart_phy_rx, soc_videosoc_uart_phy_rx_reg[7:1]};
				end
			end
		end
	end
	if (soc_videosoc_uart_phy_rx_busy) begin
		{soc_videosoc_uart_phy_uart_clk_rxen, soc_videosoc_uart_phy_phase_accumulator_rx} <= (soc_videosoc_uart_phy_phase_accumulator_rx + soc_videosoc_uart_phy_storage);
	end else begin
		{soc_videosoc_uart_phy_uart_clk_rxen, soc_videosoc_uart_phy_phase_accumulator_rx} <= 32'd2147483648;
	end
	if ((soc_videosoc_info_dna_cnt < 7'd114)) begin
		soc_videosoc_info_dna_cnt <= (soc_videosoc_info_dna_cnt + 1'd1);
		if (soc_videosoc_info_dna_cnt[0]) begin
			soc_videosoc_info_dna_status <= {soc_videosoc_info_dna_status, soc_videosoc_info_dna_do};
		end
	end
	if (soc_videosoc_info_drdy) begin
		case (soc_videosoc_info_channel)
			1'd0: begin
				soc_videosoc_info_temperature_status <= (soc_videosoc_info_data >>> 3'd4);
			end
			1'd1: begin
				soc_videosoc_info_vccint_status <= (soc_videosoc_info_data >>> 3'd4);
			end
			2'd2: begin
				soc_videosoc_info_vccaux_status <= (soc_videosoc_info_data >>> 3'd4);
			end
			3'd6: begin
				soc_videosoc_info_vccbram_status <= (soc_videosoc_info_data >>> 3'd4);
			end
		endcase
	end
	if (soc_videosoc_oled_spimaster_set_clk) begin
		soc_videosoc_oled_spi_pads_clk <= soc_videosoc_oled_spimaster_enable_cs;
	end
	if (soc_videosoc_oled_spimaster_clr_clk) begin
		soc_videosoc_oled_spi_pads_clk <= 1'd0;
		soc_videosoc_oled_spimaster_i <= 1'd0;
	end else begin
		soc_videosoc_oled_spimaster_i <= (soc_videosoc_oled_spimaster_i + 1'd1);
	end
	if (soc_videosoc_oled_spimaster_clr_cnt) begin
		soc_videosoc_oled_spimaster_cnt <= 1'd0;
	end else begin
		if (soc_videosoc_oled_spimaster_inc_cnt) begin
			soc_videosoc_oled_spimaster_cnt <= (soc_videosoc_oled_spimaster_cnt + 1'd1);
		end
	end
	if (soc_videosoc_oled_spimaster_start) begin
		soc_videosoc_oled_spimaster_sr_mosi <= soc_videosoc_oled_spimaster_mosi_storage;
	end else begin
		if ((soc_videosoc_oled_spimaster_set_clk & soc_videosoc_oled_spimaster_enable_shift)) begin
			soc_videosoc_oled_spimaster_sr_mosi <= {soc_videosoc_oled_spimaster_sr_mosi[6:0], soc_videosoc_oled_spimaster};
		end else begin
			if (soc_videosoc_oled_spimaster_clr_clk) begin
				soc_videosoc_oled_spi_pads_mosi <= soc_videosoc_oled_spimaster_sr_mosi[7];
			end
		end
	end
	vns_oled_state <= vns_oled_next_state;
	soc_videosoc_ddrphy_n_rddata_en0 <= soc_videosoc_ddrphy_dfi_p0_rddata_en;
	soc_videosoc_ddrphy_n_rddata_en1 <= soc_videosoc_ddrphy_n_rddata_en0;
	soc_videosoc_ddrphy_n_rddata_en2 <= soc_videosoc_ddrphy_n_rddata_en1;
	soc_videosoc_ddrphy_n_rddata_en3 <= soc_videosoc_ddrphy_n_rddata_en2;
	soc_videosoc_ddrphy_n_rddata_en4 <= soc_videosoc_ddrphy_n_rddata_en3;
	soc_videosoc_ddrphy_dfi_p0_rddata_valid <= soc_videosoc_ddrphy_n_rddata_en4;
	soc_videosoc_ddrphy_dfi_p1_rddata_valid <= soc_videosoc_ddrphy_n_rddata_en4;
	soc_videosoc_ddrphy_dfi_p2_rddata_valid <= soc_videosoc_ddrphy_n_rddata_en4;
	soc_videosoc_ddrphy_dfi_p3_rddata_valid <= soc_videosoc_ddrphy_n_rddata_en4;
	soc_videosoc_ddrphy_last_wrdata_en <= {soc_videosoc_ddrphy_last_wrdata_en[2:0], soc_videosoc_ddrphy_dfi_p2_wrdata_en};
	soc_videosoc_ddrphy_oe_dqs <= soc_videosoc_ddrphy_oe;
	soc_videosoc_ddrphy_oe_dq <= soc_videosoc_ddrphy_oe;
	if (soc_videosoc_sdram_inti_p0_rddata_valid) begin
		soc_videosoc_sdram_phaseinjector0_status <= soc_videosoc_sdram_inti_p0_rddata;
	end
	if (soc_videosoc_sdram_inti_p1_rddata_valid) begin
		soc_videosoc_sdram_phaseinjector1_status <= soc_videosoc_sdram_inti_p1_rddata;
	end
	if (soc_videosoc_sdram_inti_p2_rddata_valid) begin
		soc_videosoc_sdram_phaseinjector2_status <= soc_videosoc_sdram_inti_p2_rddata;
	end
	if (soc_videosoc_sdram_inti_p3_rddata_valid) begin
		soc_videosoc_sdram_phaseinjector3_status <= soc_videosoc_sdram_inti_p3_rddata;
	end
	soc_videosoc_sdram_cmd_payload_a <= 11'd1024;
	soc_videosoc_sdram_cmd_payload_ba <= 1'd0;
	soc_videosoc_sdram_cmd_payload_cas <= 1'd0;
	soc_videosoc_sdram_cmd_payload_ras <= 1'd0;
	soc_videosoc_sdram_cmd_payload_we <= 1'd0;
	soc_videosoc_sdram_seq_done <= 1'd0;
	if ((soc_videosoc_sdram_counter == 1'd1)) begin
		soc_videosoc_sdram_cmd_payload_ras <= 1'd1;
		soc_videosoc_sdram_cmd_payload_we <= 1'd1;
	end
	if ((soc_videosoc_sdram_counter == 3'd4)) begin
		soc_videosoc_sdram_cmd_payload_cas <= 1'd1;
		soc_videosoc_sdram_cmd_payload_ras <= 1'd1;
	end
	if ((soc_videosoc_sdram_counter == 5'd31)) begin
		soc_videosoc_sdram_seq_done <= 1'd1;
	end
	if ((soc_videosoc_sdram_counter != 1'd0)) begin
		soc_videosoc_sdram_counter <= (soc_videosoc_sdram_counter + 1'd1);
	end else begin
		if (soc_videosoc_sdram_seq_start) begin
			soc_videosoc_sdram_counter <= 1'd1;
		end
	end
	if (soc_videosoc_sdram_wait) begin
		if ((~soc_videosoc_sdram_done)) begin
			soc_videosoc_sdram_count <= (soc_videosoc_sdram_count - 1'd1);
		end
	end else begin
		soc_videosoc_sdram_count <= 10'd782;
	end
	vns_refresher_state <= vns_refresher_next_state;
	if (soc_videosoc_sdram_bankmachine0_track_close) begin
		soc_videosoc_sdram_bankmachine0_has_openrow <= 1'd0;
	end else begin
		if (soc_videosoc_sdram_bankmachine0_track_open) begin
			soc_videosoc_sdram_bankmachine0_has_openrow <= 1'd1;
			soc_videosoc_sdram_bankmachine0_openrow <= soc_videosoc_sdram_bankmachine0_source_payload_adr[21:7];
		end
	end
	if (((soc_videosoc_sdram_bankmachine0_syncfifo0_we & soc_videosoc_sdram_bankmachine0_syncfifo0_writable) & (~soc_videosoc_sdram_bankmachine0_replace))) begin
		soc_videosoc_sdram_bankmachine0_produce <= (soc_videosoc_sdram_bankmachine0_produce + 1'd1);
	end
	if (soc_videosoc_sdram_bankmachine0_do_read) begin
		soc_videosoc_sdram_bankmachine0_consume <= (soc_videosoc_sdram_bankmachine0_consume + 1'd1);
	end
	if (((soc_videosoc_sdram_bankmachine0_syncfifo0_we & soc_videosoc_sdram_bankmachine0_syncfifo0_writable) & (~soc_videosoc_sdram_bankmachine0_replace))) begin
		if ((~soc_videosoc_sdram_bankmachine0_do_read)) begin
			soc_videosoc_sdram_bankmachine0_level <= (soc_videosoc_sdram_bankmachine0_level + 1'd1);
		end
	end else begin
		if (soc_videosoc_sdram_bankmachine0_do_read) begin
			soc_videosoc_sdram_bankmachine0_level <= (soc_videosoc_sdram_bankmachine0_level - 1'd1);
		end
	end
	if (soc_videosoc_sdram_bankmachine0_wait) begin
		if ((~soc_videosoc_sdram_bankmachine0_done)) begin
			soc_videosoc_sdram_bankmachine0_count <= (soc_videosoc_sdram_bankmachine0_count - 1'd1);
		end
	end else begin
		soc_videosoc_sdram_bankmachine0_count <= 3'd5;
	end
	vns_bankmachine0_state <= vns_bankmachine0_next_state;
	if (soc_videosoc_sdram_bankmachine1_track_close) begin
		soc_videosoc_sdram_bankmachine1_has_openrow <= 1'd0;
	end else begin
		if (soc_videosoc_sdram_bankmachine1_track_open) begin
			soc_videosoc_sdram_bankmachine1_has_openrow <= 1'd1;
			soc_videosoc_sdram_bankmachine1_openrow <= soc_videosoc_sdram_bankmachine1_source_payload_adr[21:7];
		end
	end
	if (((soc_videosoc_sdram_bankmachine1_syncfifo1_we & soc_videosoc_sdram_bankmachine1_syncfifo1_writable) & (~soc_videosoc_sdram_bankmachine1_replace))) begin
		soc_videosoc_sdram_bankmachine1_produce <= (soc_videosoc_sdram_bankmachine1_produce + 1'd1);
	end
	if (soc_videosoc_sdram_bankmachine1_do_read) begin
		soc_videosoc_sdram_bankmachine1_consume <= (soc_videosoc_sdram_bankmachine1_consume + 1'd1);
	end
	if (((soc_videosoc_sdram_bankmachine1_syncfifo1_we & soc_videosoc_sdram_bankmachine1_syncfifo1_writable) & (~soc_videosoc_sdram_bankmachine1_replace))) begin
		if ((~soc_videosoc_sdram_bankmachine1_do_read)) begin
			soc_videosoc_sdram_bankmachine1_level <= (soc_videosoc_sdram_bankmachine1_level + 1'd1);
		end
	end else begin
		if (soc_videosoc_sdram_bankmachine1_do_read) begin
			soc_videosoc_sdram_bankmachine1_level <= (soc_videosoc_sdram_bankmachine1_level - 1'd1);
		end
	end
	if (soc_videosoc_sdram_bankmachine1_wait) begin
		if ((~soc_videosoc_sdram_bankmachine1_done)) begin
			soc_videosoc_sdram_bankmachine1_count <= (soc_videosoc_sdram_bankmachine1_count - 1'd1);
		end
	end else begin
		soc_videosoc_sdram_bankmachine1_count <= 3'd5;
	end
	vns_bankmachine1_state <= vns_bankmachine1_next_state;
	if (soc_videosoc_sdram_bankmachine2_track_close) begin
		soc_videosoc_sdram_bankmachine2_has_openrow <= 1'd0;
	end else begin
		if (soc_videosoc_sdram_bankmachine2_track_open) begin
			soc_videosoc_sdram_bankmachine2_has_openrow <= 1'd1;
			soc_videosoc_sdram_bankmachine2_openrow <= soc_videosoc_sdram_bankmachine2_source_payload_adr[21:7];
		end
	end
	if (((soc_videosoc_sdram_bankmachine2_syncfifo2_we & soc_videosoc_sdram_bankmachine2_syncfifo2_writable) & (~soc_videosoc_sdram_bankmachine2_replace))) begin
		soc_videosoc_sdram_bankmachine2_produce <= (soc_videosoc_sdram_bankmachine2_produce + 1'd1);
	end
	if (soc_videosoc_sdram_bankmachine2_do_read) begin
		soc_videosoc_sdram_bankmachine2_consume <= (soc_videosoc_sdram_bankmachine2_consume + 1'd1);
	end
	if (((soc_videosoc_sdram_bankmachine2_syncfifo2_we & soc_videosoc_sdram_bankmachine2_syncfifo2_writable) & (~soc_videosoc_sdram_bankmachine2_replace))) begin
		if ((~soc_videosoc_sdram_bankmachine2_do_read)) begin
			soc_videosoc_sdram_bankmachine2_level <= (soc_videosoc_sdram_bankmachine2_level + 1'd1);
		end
	end else begin
		if (soc_videosoc_sdram_bankmachine2_do_read) begin
			soc_videosoc_sdram_bankmachine2_level <= (soc_videosoc_sdram_bankmachine2_level - 1'd1);
		end
	end
	if (soc_videosoc_sdram_bankmachine2_wait) begin
		if ((~soc_videosoc_sdram_bankmachine2_done)) begin
			soc_videosoc_sdram_bankmachine2_count <= (soc_videosoc_sdram_bankmachine2_count - 1'd1);
		end
	end else begin
		soc_videosoc_sdram_bankmachine2_count <= 3'd5;
	end
	vns_bankmachine2_state <= vns_bankmachine2_next_state;
	if (soc_videosoc_sdram_bankmachine3_track_close) begin
		soc_videosoc_sdram_bankmachine3_has_openrow <= 1'd0;
	end else begin
		if (soc_videosoc_sdram_bankmachine3_track_open) begin
			soc_videosoc_sdram_bankmachine3_has_openrow <= 1'd1;
			soc_videosoc_sdram_bankmachine3_openrow <= soc_videosoc_sdram_bankmachine3_source_payload_adr[21:7];
		end
	end
	if (((soc_videosoc_sdram_bankmachine3_syncfifo3_we & soc_videosoc_sdram_bankmachine3_syncfifo3_writable) & (~soc_videosoc_sdram_bankmachine3_replace))) begin
		soc_videosoc_sdram_bankmachine3_produce <= (soc_videosoc_sdram_bankmachine3_produce + 1'd1);
	end
	if (soc_videosoc_sdram_bankmachine3_do_read) begin
		soc_videosoc_sdram_bankmachine3_consume <= (soc_videosoc_sdram_bankmachine3_consume + 1'd1);
	end
	if (((soc_videosoc_sdram_bankmachine3_syncfifo3_we & soc_videosoc_sdram_bankmachine3_syncfifo3_writable) & (~soc_videosoc_sdram_bankmachine3_replace))) begin
		if ((~soc_videosoc_sdram_bankmachine3_do_read)) begin
			soc_videosoc_sdram_bankmachine3_level <= (soc_videosoc_sdram_bankmachine3_level + 1'd1);
		end
	end else begin
		if (soc_videosoc_sdram_bankmachine3_do_read) begin
			soc_videosoc_sdram_bankmachine3_level <= (soc_videosoc_sdram_bankmachine3_level - 1'd1);
		end
	end
	if (soc_videosoc_sdram_bankmachine3_wait) begin
		if ((~soc_videosoc_sdram_bankmachine3_done)) begin
			soc_videosoc_sdram_bankmachine3_count <= (soc_videosoc_sdram_bankmachine3_count - 1'd1);
		end
	end else begin
		soc_videosoc_sdram_bankmachine3_count <= 3'd5;
	end
	vns_bankmachine3_state <= vns_bankmachine3_next_state;
	if (soc_videosoc_sdram_bankmachine4_track_close) begin
		soc_videosoc_sdram_bankmachine4_has_openrow <= 1'd0;
	end else begin
		if (soc_videosoc_sdram_bankmachine4_track_open) begin
			soc_videosoc_sdram_bankmachine4_has_openrow <= 1'd1;
			soc_videosoc_sdram_bankmachine4_openrow <= soc_videosoc_sdram_bankmachine4_source_payload_adr[21:7];
		end
	end
	if (((soc_videosoc_sdram_bankmachine4_syncfifo4_we & soc_videosoc_sdram_bankmachine4_syncfifo4_writable) & (~soc_videosoc_sdram_bankmachine4_replace))) begin
		soc_videosoc_sdram_bankmachine4_produce <= (soc_videosoc_sdram_bankmachine4_produce + 1'd1);
	end
	if (soc_videosoc_sdram_bankmachine4_do_read) begin
		soc_videosoc_sdram_bankmachine4_consume <= (soc_videosoc_sdram_bankmachine4_consume + 1'd1);
	end
	if (((soc_videosoc_sdram_bankmachine4_syncfifo4_we & soc_videosoc_sdram_bankmachine4_syncfifo4_writable) & (~soc_videosoc_sdram_bankmachine4_replace))) begin
		if ((~soc_videosoc_sdram_bankmachine4_do_read)) begin
			soc_videosoc_sdram_bankmachine4_level <= (soc_videosoc_sdram_bankmachine4_level + 1'd1);
		end
	end else begin
		if (soc_videosoc_sdram_bankmachine4_do_read) begin
			soc_videosoc_sdram_bankmachine4_level <= (soc_videosoc_sdram_bankmachine4_level - 1'd1);
		end
	end
	if (soc_videosoc_sdram_bankmachine4_wait) begin
		if ((~soc_videosoc_sdram_bankmachine4_done)) begin
			soc_videosoc_sdram_bankmachine4_count <= (soc_videosoc_sdram_bankmachine4_count - 1'd1);
		end
	end else begin
		soc_videosoc_sdram_bankmachine4_count <= 3'd5;
	end
	vns_bankmachine4_state <= vns_bankmachine4_next_state;
	if (soc_videosoc_sdram_bankmachine5_track_close) begin
		soc_videosoc_sdram_bankmachine5_has_openrow <= 1'd0;
	end else begin
		if (soc_videosoc_sdram_bankmachine5_track_open) begin
			soc_videosoc_sdram_bankmachine5_has_openrow <= 1'd1;
			soc_videosoc_sdram_bankmachine5_openrow <= soc_videosoc_sdram_bankmachine5_source_payload_adr[21:7];
		end
	end
	if (((soc_videosoc_sdram_bankmachine5_syncfifo5_we & soc_videosoc_sdram_bankmachine5_syncfifo5_writable) & (~soc_videosoc_sdram_bankmachine5_replace))) begin
		soc_videosoc_sdram_bankmachine5_produce <= (soc_videosoc_sdram_bankmachine5_produce + 1'd1);
	end
	if (soc_videosoc_sdram_bankmachine5_do_read) begin
		soc_videosoc_sdram_bankmachine5_consume <= (soc_videosoc_sdram_bankmachine5_consume + 1'd1);
	end
	if (((soc_videosoc_sdram_bankmachine5_syncfifo5_we & soc_videosoc_sdram_bankmachine5_syncfifo5_writable) & (~soc_videosoc_sdram_bankmachine5_replace))) begin
		if ((~soc_videosoc_sdram_bankmachine5_do_read)) begin
			soc_videosoc_sdram_bankmachine5_level <= (soc_videosoc_sdram_bankmachine5_level + 1'd1);
		end
	end else begin
		if (soc_videosoc_sdram_bankmachine5_do_read) begin
			soc_videosoc_sdram_bankmachine5_level <= (soc_videosoc_sdram_bankmachine5_level - 1'd1);
		end
	end
	if (soc_videosoc_sdram_bankmachine5_wait) begin
		if ((~soc_videosoc_sdram_bankmachine5_done)) begin
			soc_videosoc_sdram_bankmachine5_count <= (soc_videosoc_sdram_bankmachine5_count - 1'd1);
		end
	end else begin
		soc_videosoc_sdram_bankmachine5_count <= 3'd5;
	end
	vns_bankmachine5_state <= vns_bankmachine5_next_state;
	if (soc_videosoc_sdram_bankmachine6_track_close) begin
		soc_videosoc_sdram_bankmachine6_has_openrow <= 1'd0;
	end else begin
		if (soc_videosoc_sdram_bankmachine6_track_open) begin
			soc_videosoc_sdram_bankmachine6_has_openrow <= 1'd1;
			soc_videosoc_sdram_bankmachine6_openrow <= soc_videosoc_sdram_bankmachine6_source_payload_adr[21:7];
		end
	end
	if (((soc_videosoc_sdram_bankmachine6_syncfifo6_we & soc_videosoc_sdram_bankmachine6_syncfifo6_writable) & (~soc_videosoc_sdram_bankmachine6_replace))) begin
		soc_videosoc_sdram_bankmachine6_produce <= (soc_videosoc_sdram_bankmachine6_produce + 1'd1);
	end
	if (soc_videosoc_sdram_bankmachine6_do_read) begin
		soc_videosoc_sdram_bankmachine6_consume <= (soc_videosoc_sdram_bankmachine6_consume + 1'd1);
	end
	if (((soc_videosoc_sdram_bankmachine6_syncfifo6_we & soc_videosoc_sdram_bankmachine6_syncfifo6_writable) & (~soc_videosoc_sdram_bankmachine6_replace))) begin
		if ((~soc_videosoc_sdram_bankmachine6_do_read)) begin
			soc_videosoc_sdram_bankmachine6_level <= (soc_videosoc_sdram_bankmachine6_level + 1'd1);
		end
	end else begin
		if (soc_videosoc_sdram_bankmachine6_do_read) begin
			soc_videosoc_sdram_bankmachine6_level <= (soc_videosoc_sdram_bankmachine6_level - 1'd1);
		end
	end
	if (soc_videosoc_sdram_bankmachine6_wait) begin
		if ((~soc_videosoc_sdram_bankmachine6_done)) begin
			soc_videosoc_sdram_bankmachine6_count <= (soc_videosoc_sdram_bankmachine6_count - 1'd1);
		end
	end else begin
		soc_videosoc_sdram_bankmachine6_count <= 3'd5;
	end
	vns_bankmachine6_state <= vns_bankmachine6_next_state;
	if (soc_videosoc_sdram_bankmachine7_track_close) begin
		soc_videosoc_sdram_bankmachine7_has_openrow <= 1'd0;
	end else begin
		if (soc_videosoc_sdram_bankmachine7_track_open) begin
			soc_videosoc_sdram_bankmachine7_has_openrow <= 1'd1;
			soc_videosoc_sdram_bankmachine7_openrow <= soc_videosoc_sdram_bankmachine7_source_payload_adr[21:7];
		end
	end
	if (((soc_videosoc_sdram_bankmachine7_syncfifo7_we & soc_videosoc_sdram_bankmachine7_syncfifo7_writable) & (~soc_videosoc_sdram_bankmachine7_replace))) begin
		soc_videosoc_sdram_bankmachine7_produce <= (soc_videosoc_sdram_bankmachine7_produce + 1'd1);
	end
	if (soc_videosoc_sdram_bankmachine7_do_read) begin
		soc_videosoc_sdram_bankmachine7_consume <= (soc_videosoc_sdram_bankmachine7_consume + 1'd1);
	end
	if (((soc_videosoc_sdram_bankmachine7_syncfifo7_we & soc_videosoc_sdram_bankmachine7_syncfifo7_writable) & (~soc_videosoc_sdram_bankmachine7_replace))) begin
		if ((~soc_videosoc_sdram_bankmachine7_do_read)) begin
			soc_videosoc_sdram_bankmachine7_level <= (soc_videosoc_sdram_bankmachine7_level + 1'd1);
		end
	end else begin
		if (soc_videosoc_sdram_bankmachine7_do_read) begin
			soc_videosoc_sdram_bankmachine7_level <= (soc_videosoc_sdram_bankmachine7_level - 1'd1);
		end
	end
	if (soc_videosoc_sdram_bankmachine7_wait) begin
		if ((~soc_videosoc_sdram_bankmachine7_done)) begin
			soc_videosoc_sdram_bankmachine7_count <= (soc_videosoc_sdram_bankmachine7_count - 1'd1);
		end
	end else begin
		soc_videosoc_sdram_bankmachine7_count <= 3'd5;
	end
	vns_bankmachine7_state <= vns_bankmachine7_next_state;
	if ((~soc_videosoc_sdram_en0)) begin
		soc_videosoc_sdram_time0 <= 5'd31;
	end else begin
		if ((~soc_videosoc_sdram_max_time0)) begin
			soc_videosoc_sdram_time0 <= (soc_videosoc_sdram_time0 - 1'd1);
		end
	end
	if ((~soc_videosoc_sdram_en1)) begin
		soc_videosoc_sdram_time1 <= 4'd15;
	end else begin
		if ((~soc_videosoc_sdram_max_time1)) begin
			soc_videosoc_sdram_time1 <= (soc_videosoc_sdram_time1 - 1'd1);
		end
	end
	if (soc_videosoc_sdram_choose_cmd_ce) begin
		case (soc_videosoc_sdram_choose_cmd_grant)
			1'd0: begin
				if (soc_videosoc_sdram_choose_cmd_request[1]) begin
					soc_videosoc_sdram_choose_cmd_grant <= 1'd1;
				end else begin
					if (soc_videosoc_sdram_choose_cmd_request[2]) begin
						soc_videosoc_sdram_choose_cmd_grant <= 2'd2;
					end else begin
						if (soc_videosoc_sdram_choose_cmd_request[3]) begin
							soc_videosoc_sdram_choose_cmd_grant <= 2'd3;
						end else begin
							if (soc_videosoc_sdram_choose_cmd_request[4]) begin
								soc_videosoc_sdram_choose_cmd_grant <= 3'd4;
							end else begin
								if (soc_videosoc_sdram_choose_cmd_request[5]) begin
									soc_videosoc_sdram_choose_cmd_grant <= 3'd5;
								end else begin
									if (soc_videosoc_sdram_choose_cmd_request[6]) begin
										soc_videosoc_sdram_choose_cmd_grant <= 3'd6;
									end else begin
										if (soc_videosoc_sdram_choose_cmd_request[7]) begin
											soc_videosoc_sdram_choose_cmd_grant <= 3'd7;
										end
									end
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (soc_videosoc_sdram_choose_cmd_request[2]) begin
					soc_videosoc_sdram_choose_cmd_grant <= 2'd2;
				end else begin
					if (soc_videosoc_sdram_choose_cmd_request[3]) begin
						soc_videosoc_sdram_choose_cmd_grant <= 2'd3;
					end else begin
						if (soc_videosoc_sdram_choose_cmd_request[4]) begin
							soc_videosoc_sdram_choose_cmd_grant <= 3'd4;
						end else begin
							if (soc_videosoc_sdram_choose_cmd_request[5]) begin
								soc_videosoc_sdram_choose_cmd_grant <= 3'd5;
							end else begin
								if (soc_videosoc_sdram_choose_cmd_request[6]) begin
									soc_videosoc_sdram_choose_cmd_grant <= 3'd6;
								end else begin
									if (soc_videosoc_sdram_choose_cmd_request[7]) begin
										soc_videosoc_sdram_choose_cmd_grant <= 3'd7;
									end else begin
										if (soc_videosoc_sdram_choose_cmd_request[0]) begin
											soc_videosoc_sdram_choose_cmd_grant <= 1'd0;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (soc_videosoc_sdram_choose_cmd_request[3]) begin
					soc_videosoc_sdram_choose_cmd_grant <= 2'd3;
				end else begin
					if (soc_videosoc_sdram_choose_cmd_request[4]) begin
						soc_videosoc_sdram_choose_cmd_grant <= 3'd4;
					end else begin
						if (soc_videosoc_sdram_choose_cmd_request[5]) begin
							soc_videosoc_sdram_choose_cmd_grant <= 3'd5;
						end else begin
							if (soc_videosoc_sdram_choose_cmd_request[6]) begin
								soc_videosoc_sdram_choose_cmd_grant <= 3'd6;
							end else begin
								if (soc_videosoc_sdram_choose_cmd_request[7]) begin
									soc_videosoc_sdram_choose_cmd_grant <= 3'd7;
								end else begin
									if (soc_videosoc_sdram_choose_cmd_request[0]) begin
										soc_videosoc_sdram_choose_cmd_grant <= 1'd0;
									end else begin
										if (soc_videosoc_sdram_choose_cmd_request[1]) begin
											soc_videosoc_sdram_choose_cmd_grant <= 1'd1;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (soc_videosoc_sdram_choose_cmd_request[4]) begin
					soc_videosoc_sdram_choose_cmd_grant <= 3'd4;
				end else begin
					if (soc_videosoc_sdram_choose_cmd_request[5]) begin
						soc_videosoc_sdram_choose_cmd_grant <= 3'd5;
					end else begin
						if (soc_videosoc_sdram_choose_cmd_request[6]) begin
							soc_videosoc_sdram_choose_cmd_grant <= 3'd6;
						end else begin
							if (soc_videosoc_sdram_choose_cmd_request[7]) begin
								soc_videosoc_sdram_choose_cmd_grant <= 3'd7;
							end else begin
								if (soc_videosoc_sdram_choose_cmd_request[0]) begin
									soc_videosoc_sdram_choose_cmd_grant <= 1'd0;
								end else begin
									if (soc_videosoc_sdram_choose_cmd_request[1]) begin
										soc_videosoc_sdram_choose_cmd_grant <= 1'd1;
									end else begin
										if (soc_videosoc_sdram_choose_cmd_request[2]) begin
											soc_videosoc_sdram_choose_cmd_grant <= 2'd2;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (soc_videosoc_sdram_choose_cmd_request[5]) begin
					soc_videosoc_sdram_choose_cmd_grant <= 3'd5;
				end else begin
					if (soc_videosoc_sdram_choose_cmd_request[6]) begin
						soc_videosoc_sdram_choose_cmd_grant <= 3'd6;
					end else begin
						if (soc_videosoc_sdram_choose_cmd_request[7]) begin
							soc_videosoc_sdram_choose_cmd_grant <= 3'd7;
						end else begin
							if (soc_videosoc_sdram_choose_cmd_request[0]) begin
								soc_videosoc_sdram_choose_cmd_grant <= 1'd0;
							end else begin
								if (soc_videosoc_sdram_choose_cmd_request[1]) begin
									soc_videosoc_sdram_choose_cmd_grant <= 1'd1;
								end else begin
									if (soc_videosoc_sdram_choose_cmd_request[2]) begin
										soc_videosoc_sdram_choose_cmd_grant <= 2'd2;
									end else begin
										if (soc_videosoc_sdram_choose_cmd_request[3]) begin
											soc_videosoc_sdram_choose_cmd_grant <= 2'd3;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (soc_videosoc_sdram_choose_cmd_request[6]) begin
					soc_videosoc_sdram_choose_cmd_grant <= 3'd6;
				end else begin
					if (soc_videosoc_sdram_choose_cmd_request[7]) begin
						soc_videosoc_sdram_choose_cmd_grant <= 3'd7;
					end else begin
						if (soc_videosoc_sdram_choose_cmd_request[0]) begin
							soc_videosoc_sdram_choose_cmd_grant <= 1'd0;
						end else begin
							if (soc_videosoc_sdram_choose_cmd_request[1]) begin
								soc_videosoc_sdram_choose_cmd_grant <= 1'd1;
							end else begin
								if (soc_videosoc_sdram_choose_cmd_request[2]) begin
									soc_videosoc_sdram_choose_cmd_grant <= 2'd2;
								end else begin
									if (soc_videosoc_sdram_choose_cmd_request[3]) begin
										soc_videosoc_sdram_choose_cmd_grant <= 2'd3;
									end else begin
										if (soc_videosoc_sdram_choose_cmd_request[4]) begin
											soc_videosoc_sdram_choose_cmd_grant <= 3'd4;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd6: begin
				if (soc_videosoc_sdram_choose_cmd_request[7]) begin
					soc_videosoc_sdram_choose_cmd_grant <= 3'd7;
				end else begin
					if (soc_videosoc_sdram_choose_cmd_request[0]) begin
						soc_videosoc_sdram_choose_cmd_grant <= 1'd0;
					end else begin
						if (soc_videosoc_sdram_choose_cmd_request[1]) begin
							soc_videosoc_sdram_choose_cmd_grant <= 1'd1;
						end else begin
							if (soc_videosoc_sdram_choose_cmd_request[2]) begin
								soc_videosoc_sdram_choose_cmd_grant <= 2'd2;
							end else begin
								if (soc_videosoc_sdram_choose_cmd_request[3]) begin
									soc_videosoc_sdram_choose_cmd_grant <= 2'd3;
								end else begin
									if (soc_videosoc_sdram_choose_cmd_request[4]) begin
										soc_videosoc_sdram_choose_cmd_grant <= 3'd4;
									end else begin
										if (soc_videosoc_sdram_choose_cmd_request[5]) begin
											soc_videosoc_sdram_choose_cmd_grant <= 3'd5;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd7: begin
				if (soc_videosoc_sdram_choose_cmd_request[0]) begin
					soc_videosoc_sdram_choose_cmd_grant <= 1'd0;
				end else begin
					if (soc_videosoc_sdram_choose_cmd_request[1]) begin
						soc_videosoc_sdram_choose_cmd_grant <= 1'd1;
					end else begin
						if (soc_videosoc_sdram_choose_cmd_request[2]) begin
							soc_videosoc_sdram_choose_cmd_grant <= 2'd2;
						end else begin
							if (soc_videosoc_sdram_choose_cmd_request[3]) begin
								soc_videosoc_sdram_choose_cmd_grant <= 2'd3;
							end else begin
								if (soc_videosoc_sdram_choose_cmd_request[4]) begin
									soc_videosoc_sdram_choose_cmd_grant <= 3'd4;
								end else begin
									if (soc_videosoc_sdram_choose_cmd_request[5]) begin
										soc_videosoc_sdram_choose_cmd_grant <= 3'd5;
									end else begin
										if (soc_videosoc_sdram_choose_cmd_request[6]) begin
											soc_videosoc_sdram_choose_cmd_grant <= 3'd6;
										end
									end
								end
							end
						end
					end
				end
			end
		endcase
	end
	if (soc_videosoc_sdram_choose_req_ce) begin
		case (soc_videosoc_sdram_choose_req_grant)
			1'd0: begin
				if (soc_videosoc_sdram_choose_req_request[1]) begin
					soc_videosoc_sdram_choose_req_grant <= 1'd1;
				end else begin
					if (soc_videosoc_sdram_choose_req_request[2]) begin
						soc_videosoc_sdram_choose_req_grant <= 2'd2;
					end else begin
						if (soc_videosoc_sdram_choose_req_request[3]) begin
							soc_videosoc_sdram_choose_req_grant <= 2'd3;
						end else begin
							if (soc_videosoc_sdram_choose_req_request[4]) begin
								soc_videosoc_sdram_choose_req_grant <= 3'd4;
							end else begin
								if (soc_videosoc_sdram_choose_req_request[5]) begin
									soc_videosoc_sdram_choose_req_grant <= 3'd5;
								end else begin
									if (soc_videosoc_sdram_choose_req_request[6]) begin
										soc_videosoc_sdram_choose_req_grant <= 3'd6;
									end else begin
										if (soc_videosoc_sdram_choose_req_request[7]) begin
											soc_videosoc_sdram_choose_req_grant <= 3'd7;
										end
									end
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (soc_videosoc_sdram_choose_req_request[2]) begin
					soc_videosoc_sdram_choose_req_grant <= 2'd2;
				end else begin
					if (soc_videosoc_sdram_choose_req_request[3]) begin
						soc_videosoc_sdram_choose_req_grant <= 2'd3;
					end else begin
						if (soc_videosoc_sdram_choose_req_request[4]) begin
							soc_videosoc_sdram_choose_req_grant <= 3'd4;
						end else begin
							if (soc_videosoc_sdram_choose_req_request[5]) begin
								soc_videosoc_sdram_choose_req_grant <= 3'd5;
							end else begin
								if (soc_videosoc_sdram_choose_req_request[6]) begin
									soc_videosoc_sdram_choose_req_grant <= 3'd6;
								end else begin
									if (soc_videosoc_sdram_choose_req_request[7]) begin
										soc_videosoc_sdram_choose_req_grant <= 3'd7;
									end else begin
										if (soc_videosoc_sdram_choose_req_request[0]) begin
											soc_videosoc_sdram_choose_req_grant <= 1'd0;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (soc_videosoc_sdram_choose_req_request[3]) begin
					soc_videosoc_sdram_choose_req_grant <= 2'd3;
				end else begin
					if (soc_videosoc_sdram_choose_req_request[4]) begin
						soc_videosoc_sdram_choose_req_grant <= 3'd4;
					end else begin
						if (soc_videosoc_sdram_choose_req_request[5]) begin
							soc_videosoc_sdram_choose_req_grant <= 3'd5;
						end else begin
							if (soc_videosoc_sdram_choose_req_request[6]) begin
								soc_videosoc_sdram_choose_req_grant <= 3'd6;
							end else begin
								if (soc_videosoc_sdram_choose_req_request[7]) begin
									soc_videosoc_sdram_choose_req_grant <= 3'd7;
								end else begin
									if (soc_videosoc_sdram_choose_req_request[0]) begin
										soc_videosoc_sdram_choose_req_grant <= 1'd0;
									end else begin
										if (soc_videosoc_sdram_choose_req_request[1]) begin
											soc_videosoc_sdram_choose_req_grant <= 1'd1;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (soc_videosoc_sdram_choose_req_request[4]) begin
					soc_videosoc_sdram_choose_req_grant <= 3'd4;
				end else begin
					if (soc_videosoc_sdram_choose_req_request[5]) begin
						soc_videosoc_sdram_choose_req_grant <= 3'd5;
					end else begin
						if (soc_videosoc_sdram_choose_req_request[6]) begin
							soc_videosoc_sdram_choose_req_grant <= 3'd6;
						end else begin
							if (soc_videosoc_sdram_choose_req_request[7]) begin
								soc_videosoc_sdram_choose_req_grant <= 3'd7;
							end else begin
								if (soc_videosoc_sdram_choose_req_request[0]) begin
									soc_videosoc_sdram_choose_req_grant <= 1'd0;
								end else begin
									if (soc_videosoc_sdram_choose_req_request[1]) begin
										soc_videosoc_sdram_choose_req_grant <= 1'd1;
									end else begin
										if (soc_videosoc_sdram_choose_req_request[2]) begin
											soc_videosoc_sdram_choose_req_grant <= 2'd2;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (soc_videosoc_sdram_choose_req_request[5]) begin
					soc_videosoc_sdram_choose_req_grant <= 3'd5;
				end else begin
					if (soc_videosoc_sdram_choose_req_request[6]) begin
						soc_videosoc_sdram_choose_req_grant <= 3'd6;
					end else begin
						if (soc_videosoc_sdram_choose_req_request[7]) begin
							soc_videosoc_sdram_choose_req_grant <= 3'd7;
						end else begin
							if (soc_videosoc_sdram_choose_req_request[0]) begin
								soc_videosoc_sdram_choose_req_grant <= 1'd0;
							end else begin
								if (soc_videosoc_sdram_choose_req_request[1]) begin
									soc_videosoc_sdram_choose_req_grant <= 1'd1;
								end else begin
									if (soc_videosoc_sdram_choose_req_request[2]) begin
										soc_videosoc_sdram_choose_req_grant <= 2'd2;
									end else begin
										if (soc_videosoc_sdram_choose_req_request[3]) begin
											soc_videosoc_sdram_choose_req_grant <= 2'd3;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (soc_videosoc_sdram_choose_req_request[6]) begin
					soc_videosoc_sdram_choose_req_grant <= 3'd6;
				end else begin
					if (soc_videosoc_sdram_choose_req_request[7]) begin
						soc_videosoc_sdram_choose_req_grant <= 3'd7;
					end else begin
						if (soc_videosoc_sdram_choose_req_request[0]) begin
							soc_videosoc_sdram_choose_req_grant <= 1'd0;
						end else begin
							if (soc_videosoc_sdram_choose_req_request[1]) begin
								soc_videosoc_sdram_choose_req_grant <= 1'd1;
							end else begin
								if (soc_videosoc_sdram_choose_req_request[2]) begin
									soc_videosoc_sdram_choose_req_grant <= 2'd2;
								end else begin
									if (soc_videosoc_sdram_choose_req_request[3]) begin
										soc_videosoc_sdram_choose_req_grant <= 2'd3;
									end else begin
										if (soc_videosoc_sdram_choose_req_request[4]) begin
											soc_videosoc_sdram_choose_req_grant <= 3'd4;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd6: begin
				if (soc_videosoc_sdram_choose_req_request[7]) begin
					soc_videosoc_sdram_choose_req_grant <= 3'd7;
				end else begin
					if (soc_videosoc_sdram_choose_req_request[0]) begin
						soc_videosoc_sdram_choose_req_grant <= 1'd0;
					end else begin
						if (soc_videosoc_sdram_choose_req_request[1]) begin
							soc_videosoc_sdram_choose_req_grant <= 1'd1;
						end else begin
							if (soc_videosoc_sdram_choose_req_request[2]) begin
								soc_videosoc_sdram_choose_req_grant <= 2'd2;
							end else begin
								if (soc_videosoc_sdram_choose_req_request[3]) begin
									soc_videosoc_sdram_choose_req_grant <= 2'd3;
								end else begin
									if (soc_videosoc_sdram_choose_req_request[4]) begin
										soc_videosoc_sdram_choose_req_grant <= 3'd4;
									end else begin
										if (soc_videosoc_sdram_choose_req_request[5]) begin
											soc_videosoc_sdram_choose_req_grant <= 3'd5;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd7: begin
				if (soc_videosoc_sdram_choose_req_request[0]) begin
					soc_videosoc_sdram_choose_req_grant <= 1'd0;
				end else begin
					if (soc_videosoc_sdram_choose_req_request[1]) begin
						soc_videosoc_sdram_choose_req_grant <= 1'd1;
					end else begin
						if (soc_videosoc_sdram_choose_req_request[2]) begin
							soc_videosoc_sdram_choose_req_grant <= 2'd2;
						end else begin
							if (soc_videosoc_sdram_choose_req_request[3]) begin
								soc_videosoc_sdram_choose_req_grant <= 2'd3;
							end else begin
								if (soc_videosoc_sdram_choose_req_request[4]) begin
									soc_videosoc_sdram_choose_req_grant <= 3'd4;
								end else begin
									if (soc_videosoc_sdram_choose_req_request[5]) begin
										soc_videosoc_sdram_choose_req_grant <= 3'd5;
									end else begin
										if (soc_videosoc_sdram_choose_req_request[6]) begin
											soc_videosoc_sdram_choose_req_grant <= 3'd6;
										end
									end
								end
							end
						end
					end
				end
			end
		endcase
	end
	soc_videosoc_sdram_dfi_p0_address <= vns_sync_rhs_array_muxed0;
	soc_videosoc_sdram_dfi_p0_bank <= vns_sync_rhs_array_muxed1;
	soc_videosoc_sdram_dfi_p0_cas_n <= (~vns_sync_rhs_array_muxed2);
	soc_videosoc_sdram_dfi_p0_ras_n <= (~vns_sync_rhs_array_muxed3);
	soc_videosoc_sdram_dfi_p0_we_n <= (~vns_sync_rhs_array_muxed4);
	soc_videosoc_sdram_dfi_p0_rddata_en <= vns_sync_rhs_array_muxed5;
	soc_videosoc_sdram_dfi_p0_wrdata_en <= vns_sync_rhs_array_muxed6;
	soc_videosoc_sdram_dfi_p1_address <= vns_sync_rhs_array_muxed7;
	soc_videosoc_sdram_dfi_p1_bank <= vns_sync_rhs_array_muxed8;
	soc_videosoc_sdram_dfi_p1_cas_n <= (~vns_sync_rhs_array_muxed9);
	soc_videosoc_sdram_dfi_p1_ras_n <= (~vns_sync_rhs_array_muxed10);
	soc_videosoc_sdram_dfi_p1_we_n <= (~vns_sync_rhs_array_muxed11);
	soc_videosoc_sdram_dfi_p1_rddata_en <= vns_sync_rhs_array_muxed12;
	soc_videosoc_sdram_dfi_p1_wrdata_en <= vns_sync_rhs_array_muxed13;
	soc_videosoc_sdram_dfi_p2_address <= vns_sync_rhs_array_muxed14;
	soc_videosoc_sdram_dfi_p2_bank <= vns_sync_rhs_array_muxed15;
	soc_videosoc_sdram_dfi_p2_cas_n <= (~vns_sync_rhs_array_muxed16);
	soc_videosoc_sdram_dfi_p2_ras_n <= (~vns_sync_rhs_array_muxed17);
	soc_videosoc_sdram_dfi_p2_we_n <= (~vns_sync_rhs_array_muxed18);
	soc_videosoc_sdram_dfi_p2_rddata_en <= vns_sync_rhs_array_muxed19;
	soc_videosoc_sdram_dfi_p2_wrdata_en <= vns_sync_rhs_array_muxed20;
	soc_videosoc_sdram_dfi_p3_address <= vns_sync_rhs_array_muxed21;
	soc_videosoc_sdram_dfi_p3_bank <= vns_sync_rhs_array_muxed22;
	soc_videosoc_sdram_dfi_p3_cas_n <= (~vns_sync_rhs_array_muxed23);
	soc_videosoc_sdram_dfi_p3_ras_n <= (~vns_sync_rhs_array_muxed24);
	soc_videosoc_sdram_dfi_p3_we_n <= (~vns_sync_rhs_array_muxed25);
	soc_videosoc_sdram_dfi_p3_rddata_en <= vns_sync_rhs_array_muxed26;
	soc_videosoc_sdram_dfi_p3_wrdata_en <= vns_sync_rhs_array_muxed27;
	vns_multiplexer_state <= vns_multiplexer_next_state;
	soc_videosoc_sdram_bandwidth_cmd_valid <= soc_videosoc_sdram_choose_req_cmd_valid;
	soc_videosoc_sdram_bandwidth_cmd_ready <= soc_videosoc_sdram_choose_req_cmd_ready;
	soc_videosoc_sdram_bandwidth_cmd_is_read <= soc_videosoc_sdram_choose_req_cmd_payload_is_read;
	soc_videosoc_sdram_bandwidth_cmd_is_write <= soc_videosoc_sdram_choose_req_cmd_payload_is_write;
	{soc_videosoc_sdram_bandwidth_period, soc_videosoc_sdram_bandwidth_counter} <= (soc_videosoc_sdram_bandwidth_counter + 1'd1);
	if (soc_videosoc_sdram_bandwidth_period) begin
		soc_videosoc_sdram_bandwidth_nreads_r <= soc_videosoc_sdram_bandwidth_nreads;
		soc_videosoc_sdram_bandwidth_nwrites_r <= soc_videosoc_sdram_bandwidth_nwrites;
		soc_videosoc_sdram_bandwidth_nreads <= 1'd0;
		soc_videosoc_sdram_bandwidth_nwrites <= 1'd0;
	end else begin
		if ((soc_videosoc_sdram_bandwidth_cmd_valid & soc_videosoc_sdram_bandwidth_cmd_ready)) begin
			if (soc_videosoc_sdram_bandwidth_cmd_is_read) begin
				soc_videosoc_sdram_bandwidth_nreads <= (soc_videosoc_sdram_bandwidth_nreads + 1'd1);
			end
			if (soc_videosoc_sdram_bandwidth_cmd_is_write) begin
				soc_videosoc_sdram_bandwidth_nwrites <= (soc_videosoc_sdram_bandwidth_nwrites + 1'd1);
			end
		end
	end
	if (soc_videosoc_sdram_bandwidth_update_re) begin
		soc_videosoc_sdram_bandwidth_nreads_status <= soc_videosoc_sdram_bandwidth_nreads_r;
		soc_videosoc_sdram_bandwidth_nwrites_status <= soc_videosoc_sdram_bandwidth_nwrites_r;
	end
	vns_new_master_wdata_ready0 <= ((((((((1'd0 | ((vns_roundrobin0_grant == 1'd0) & soc_videosoc_sdram_interface_bank0_wdata_ready)) | ((vns_roundrobin1_grant == 1'd0) & soc_videosoc_sdram_interface_bank1_wdata_ready)) | ((vns_roundrobin2_grant == 1'd0) & soc_videosoc_sdram_interface_bank2_wdata_ready)) | ((vns_roundrobin3_grant == 1'd0) & soc_videosoc_sdram_interface_bank3_wdata_ready)) | ((vns_roundrobin4_grant == 1'd0) & soc_videosoc_sdram_interface_bank4_wdata_ready)) | ((vns_roundrobin5_grant == 1'd0) & soc_videosoc_sdram_interface_bank5_wdata_ready)) | ((vns_roundrobin6_grant == 1'd0) & soc_videosoc_sdram_interface_bank6_wdata_ready)) | ((vns_roundrobin7_grant == 1'd0) & soc_videosoc_sdram_interface_bank7_wdata_ready));
	vns_new_master_wdata_ready1 <= vns_new_master_wdata_ready0;
	vns_new_master_wdata_ready2 <= vns_new_master_wdata_ready1;
	vns_new_master_wdata_ready3 <= ((((((((1'd0 | ((vns_roundrobin0_grant == 1'd1) & soc_videosoc_sdram_interface_bank0_wdata_ready)) | ((vns_roundrobin1_grant == 1'd1) & soc_videosoc_sdram_interface_bank1_wdata_ready)) | ((vns_roundrobin2_grant == 1'd1) & soc_videosoc_sdram_interface_bank2_wdata_ready)) | ((vns_roundrobin3_grant == 1'd1) & soc_videosoc_sdram_interface_bank3_wdata_ready)) | ((vns_roundrobin4_grant == 1'd1) & soc_videosoc_sdram_interface_bank4_wdata_ready)) | ((vns_roundrobin5_grant == 1'd1) & soc_videosoc_sdram_interface_bank5_wdata_ready)) | ((vns_roundrobin6_grant == 1'd1) & soc_videosoc_sdram_interface_bank6_wdata_ready)) | ((vns_roundrobin7_grant == 1'd1) & soc_videosoc_sdram_interface_bank7_wdata_ready));
	vns_new_master_wdata_ready4 <= vns_new_master_wdata_ready3;
	vns_new_master_wdata_ready5 <= vns_new_master_wdata_ready4;
	vns_new_master_wdata_ready6 <= ((((((((1'd0 | ((vns_roundrobin0_grant == 2'd2) & soc_videosoc_sdram_interface_bank0_wdata_ready)) | ((vns_roundrobin1_grant == 2'd2) & soc_videosoc_sdram_interface_bank1_wdata_ready)) | ((vns_roundrobin2_grant == 2'd2) & soc_videosoc_sdram_interface_bank2_wdata_ready)) | ((vns_roundrobin3_grant == 2'd2) & soc_videosoc_sdram_interface_bank3_wdata_ready)) | ((vns_roundrobin4_grant == 2'd2) & soc_videosoc_sdram_interface_bank4_wdata_ready)) | ((vns_roundrobin5_grant == 2'd2) & soc_videosoc_sdram_interface_bank5_wdata_ready)) | ((vns_roundrobin6_grant == 2'd2) & soc_videosoc_sdram_interface_bank6_wdata_ready)) | ((vns_roundrobin7_grant == 2'd2) & soc_videosoc_sdram_interface_bank7_wdata_ready));
	vns_new_master_wdata_ready7 <= vns_new_master_wdata_ready6;
	vns_new_master_wdata_ready8 <= vns_new_master_wdata_ready7;
	vns_new_master_rdata_valid0 <= ((((((((1'd0 | ((vns_roundrobin0_grant == 1'd0) & soc_videosoc_sdram_interface_bank0_rdata_valid)) | ((vns_roundrobin1_grant == 1'd0) & soc_videosoc_sdram_interface_bank1_rdata_valid)) | ((vns_roundrobin2_grant == 1'd0) & soc_videosoc_sdram_interface_bank2_rdata_valid)) | ((vns_roundrobin3_grant == 1'd0) & soc_videosoc_sdram_interface_bank3_rdata_valid)) | ((vns_roundrobin4_grant == 1'd0) & soc_videosoc_sdram_interface_bank4_rdata_valid)) | ((vns_roundrobin5_grant == 1'd0) & soc_videosoc_sdram_interface_bank5_rdata_valid)) | ((vns_roundrobin6_grant == 1'd0) & soc_videosoc_sdram_interface_bank6_rdata_valid)) | ((vns_roundrobin7_grant == 1'd0) & soc_videosoc_sdram_interface_bank7_rdata_valid));
	vns_new_master_rdata_valid1 <= vns_new_master_rdata_valid0;
	vns_new_master_rdata_valid2 <= vns_new_master_rdata_valid1;
	vns_new_master_rdata_valid3 <= vns_new_master_rdata_valid2;
	vns_new_master_rdata_valid4 <= vns_new_master_rdata_valid3;
	vns_new_master_rdata_valid5 <= vns_new_master_rdata_valid4;
	vns_new_master_rdata_valid6 <= vns_new_master_rdata_valid5;
	vns_new_master_rdata_valid7 <= ((((((((1'd0 | ((vns_roundrobin0_grant == 1'd1) & soc_videosoc_sdram_interface_bank0_rdata_valid)) | ((vns_roundrobin1_grant == 1'd1) & soc_videosoc_sdram_interface_bank1_rdata_valid)) | ((vns_roundrobin2_grant == 1'd1) & soc_videosoc_sdram_interface_bank2_rdata_valid)) | ((vns_roundrobin3_grant == 1'd1) & soc_videosoc_sdram_interface_bank3_rdata_valid)) | ((vns_roundrobin4_grant == 1'd1) & soc_videosoc_sdram_interface_bank4_rdata_valid)) | ((vns_roundrobin5_grant == 1'd1) & soc_videosoc_sdram_interface_bank5_rdata_valid)) | ((vns_roundrobin6_grant == 1'd1) & soc_videosoc_sdram_interface_bank6_rdata_valid)) | ((vns_roundrobin7_grant == 1'd1) & soc_videosoc_sdram_interface_bank7_rdata_valid));
	vns_new_master_rdata_valid8 <= vns_new_master_rdata_valid7;
	vns_new_master_rdata_valid9 <= vns_new_master_rdata_valid8;
	vns_new_master_rdata_valid10 <= vns_new_master_rdata_valid9;
	vns_new_master_rdata_valid11 <= vns_new_master_rdata_valid10;
	vns_new_master_rdata_valid12 <= vns_new_master_rdata_valid11;
	vns_new_master_rdata_valid13 <= vns_new_master_rdata_valid12;
	vns_new_master_rdata_valid14 <= ((((((((1'd0 | ((vns_roundrobin0_grant == 2'd2) & soc_videosoc_sdram_interface_bank0_rdata_valid)) | ((vns_roundrobin1_grant == 2'd2) & soc_videosoc_sdram_interface_bank1_rdata_valid)) | ((vns_roundrobin2_grant == 2'd2) & soc_videosoc_sdram_interface_bank2_rdata_valid)) | ((vns_roundrobin3_grant == 2'd2) & soc_videosoc_sdram_interface_bank3_rdata_valid)) | ((vns_roundrobin4_grant == 2'd2) & soc_videosoc_sdram_interface_bank4_rdata_valid)) | ((vns_roundrobin5_grant == 2'd2) & soc_videosoc_sdram_interface_bank5_rdata_valid)) | ((vns_roundrobin6_grant == 2'd2) & soc_videosoc_sdram_interface_bank6_rdata_valid)) | ((vns_roundrobin7_grant == 2'd2) & soc_videosoc_sdram_interface_bank7_rdata_valid));
	vns_new_master_rdata_valid15 <= vns_new_master_rdata_valid14;
	vns_new_master_rdata_valid16 <= vns_new_master_rdata_valid15;
	vns_new_master_rdata_valid17 <= vns_new_master_rdata_valid16;
	vns_new_master_rdata_valid18 <= vns_new_master_rdata_valid17;
	vns_new_master_rdata_valid19 <= vns_new_master_rdata_valid18;
	vns_new_master_rdata_valid20 <= vns_new_master_rdata_valid19;
	soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_binary <= soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next_binary;
	soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q <= soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_next;
	soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_binary <= soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next_binary;
	soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q <= soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_next;
	if (vns_roundrobin0_ce) begin
		case (vns_roundrobin0_grant)
			1'd0: begin
				if (vns_roundrobin0_request[1]) begin
					vns_roundrobin0_grant <= 1'd1;
				end else begin
					if (vns_roundrobin0_request[2]) begin
						vns_roundrobin0_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin0_request[2]) begin
					vns_roundrobin0_grant <= 2'd2;
				end else begin
					if (vns_roundrobin0_request[0]) begin
						vns_roundrobin0_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin0_request[0]) begin
					vns_roundrobin0_grant <= 1'd0;
				end else begin
					if (vns_roundrobin0_request[1]) begin
						vns_roundrobin0_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (vns_roundrobin1_ce) begin
		case (vns_roundrobin1_grant)
			1'd0: begin
				if (vns_roundrobin1_request[1]) begin
					vns_roundrobin1_grant <= 1'd1;
				end else begin
					if (vns_roundrobin1_request[2]) begin
						vns_roundrobin1_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin1_request[2]) begin
					vns_roundrobin1_grant <= 2'd2;
				end else begin
					if (vns_roundrobin1_request[0]) begin
						vns_roundrobin1_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin1_request[0]) begin
					vns_roundrobin1_grant <= 1'd0;
				end else begin
					if (vns_roundrobin1_request[1]) begin
						vns_roundrobin1_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (vns_roundrobin2_ce) begin
		case (vns_roundrobin2_grant)
			1'd0: begin
				if (vns_roundrobin2_request[1]) begin
					vns_roundrobin2_grant <= 1'd1;
				end else begin
					if (vns_roundrobin2_request[2]) begin
						vns_roundrobin2_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin2_request[2]) begin
					vns_roundrobin2_grant <= 2'd2;
				end else begin
					if (vns_roundrobin2_request[0]) begin
						vns_roundrobin2_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin2_request[0]) begin
					vns_roundrobin2_grant <= 1'd0;
				end else begin
					if (vns_roundrobin2_request[1]) begin
						vns_roundrobin2_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (vns_roundrobin3_ce) begin
		case (vns_roundrobin3_grant)
			1'd0: begin
				if (vns_roundrobin3_request[1]) begin
					vns_roundrobin3_grant <= 1'd1;
				end else begin
					if (vns_roundrobin3_request[2]) begin
						vns_roundrobin3_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin3_request[2]) begin
					vns_roundrobin3_grant <= 2'd2;
				end else begin
					if (vns_roundrobin3_request[0]) begin
						vns_roundrobin3_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin3_request[0]) begin
					vns_roundrobin3_grant <= 1'd0;
				end else begin
					if (vns_roundrobin3_request[1]) begin
						vns_roundrobin3_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (vns_roundrobin4_ce) begin
		case (vns_roundrobin4_grant)
			1'd0: begin
				if (vns_roundrobin4_request[1]) begin
					vns_roundrobin4_grant <= 1'd1;
				end else begin
					if (vns_roundrobin4_request[2]) begin
						vns_roundrobin4_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin4_request[2]) begin
					vns_roundrobin4_grant <= 2'd2;
				end else begin
					if (vns_roundrobin4_request[0]) begin
						vns_roundrobin4_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin4_request[0]) begin
					vns_roundrobin4_grant <= 1'd0;
				end else begin
					if (vns_roundrobin4_request[1]) begin
						vns_roundrobin4_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (vns_roundrobin5_ce) begin
		case (vns_roundrobin5_grant)
			1'd0: begin
				if (vns_roundrobin5_request[1]) begin
					vns_roundrobin5_grant <= 1'd1;
				end else begin
					if (vns_roundrobin5_request[2]) begin
						vns_roundrobin5_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin5_request[2]) begin
					vns_roundrobin5_grant <= 2'd2;
				end else begin
					if (vns_roundrobin5_request[0]) begin
						vns_roundrobin5_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin5_request[0]) begin
					vns_roundrobin5_grant <= 1'd0;
				end else begin
					if (vns_roundrobin5_request[1]) begin
						vns_roundrobin5_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (vns_roundrobin6_ce) begin
		case (vns_roundrobin6_grant)
			1'd0: begin
				if (vns_roundrobin6_request[1]) begin
					vns_roundrobin6_grant <= 1'd1;
				end else begin
					if (vns_roundrobin6_request[2]) begin
						vns_roundrobin6_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin6_request[2]) begin
					vns_roundrobin6_grant <= 2'd2;
				end else begin
					if (vns_roundrobin6_request[0]) begin
						vns_roundrobin6_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin6_request[0]) begin
					vns_roundrobin6_grant <= 1'd0;
				end else begin
					if (vns_roundrobin6_request[1]) begin
						vns_roundrobin6_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	if (vns_roundrobin7_ce) begin
		case (vns_roundrobin7_grant)
			1'd0: begin
				if (vns_roundrobin7_request[1]) begin
					vns_roundrobin7_grant <= 1'd1;
				end else begin
					if (vns_roundrobin7_request[2]) begin
						vns_roundrobin7_grant <= 2'd2;
					end
				end
			end
			1'd1: begin
				if (vns_roundrobin7_request[2]) begin
					vns_roundrobin7_grant <= 2'd2;
				end else begin
					if (vns_roundrobin7_request[0]) begin
						vns_roundrobin7_grant <= 1'd0;
					end
				end
			end
			2'd2: begin
				if (vns_roundrobin7_request[0]) begin
					vns_roundrobin7_grant <= 1'd0;
				end else begin
					if (vns_roundrobin7_request[1]) begin
						vns_roundrobin7_grant <= 1'd1;
					end
				end
			end
		endcase
	end
	soc_videosoc_adr_offset_r <= soc_videosoc_interface0_wb_sdram_adr[1:0];
	vns_fullmemorywe_state <= vns_fullmemorywe_next_state;
	vns_litedramwishbonebridge_state <= vns_litedramwishbonebridge_next_state;
	if ((soc_videosoc_i == 1'd0)) begin
		soc_videosoc_clk1 <= 1'd1;
		soc_videosoc_miso <= spiflash_1x_miso;
	end
	if ((soc_videosoc_i == 1'd1)) begin
		soc_videosoc_i <= 1'd0;
		soc_videosoc_clk1 <= 1'd0;
		soc_videosoc_sr <= {soc_videosoc_sr[30:0], soc_videosoc_miso};
	end else begin
		soc_videosoc_i <= (soc_videosoc_i + 1'd1);
	end
	if ((((soc_videosoc_bus_cyc & soc_videosoc_bus_stb) & (soc_videosoc_i == 1'd1)) & (soc_videosoc_counter == 1'd0))) begin
		soc_videosoc_cs_n <= 1'd0;
		soc_videosoc_sr[31:24] <= 4'd11;
	end
	if ((soc_videosoc_counter == 5'd16)) begin
		soc_videosoc_sr[31:8] <= {soc_videosoc_bus_adr, {2{1'd0}}};
	end
	if ((soc_videosoc_counter == 7'd64)) begin
	end
	if ((soc_videosoc_counter == 8'd146)) begin
		soc_videosoc_bus_ack <= 1'd1;
		soc_videosoc_cs_n <= 1'd1;
	end
	if ((soc_videosoc_counter == 8'd147)) begin
		soc_videosoc_bus_ack <= 1'd0;
	end
	if ((soc_videosoc_counter == 8'd149)) begin
	end
	if ((soc_videosoc_counter == 8'd149)) begin
		soc_videosoc_counter <= 1'd0;
	end else begin
		if ((soc_videosoc_counter != 1'd0)) begin
			soc_videosoc_counter <= (soc_videosoc_counter + 1'd1);
		end else begin
			if (((soc_videosoc_bus_cyc & soc_videosoc_bus_stb) & (soc_videosoc_i == 1'd1))) begin
				soc_videosoc_counter <= 1'd1;
			end
		end
	end
	if (soc_ethphy_counter_ce) begin
		soc_ethphy_counter <= (soc_ethphy_counter + 1'd1);
	end
	soc_ethmac_tx_cdc_graycounter0_q_binary <= soc_ethmac_tx_cdc_graycounter0_q_next_binary;
	soc_ethmac_tx_cdc_graycounter0_q <= soc_ethmac_tx_cdc_graycounter0_q_next;
	soc_ethmac_rx_cdc_graycounter1_q_binary <= soc_ethmac_rx_cdc_graycounter1_q_next_binary;
	soc_ethmac_rx_cdc_graycounter1_q <= soc_ethmac_rx_cdc_graycounter1_q_next;
	if (soc_ethmac_writer_counter_reset) begin
		soc_ethmac_writer_counter <= 1'd0;
	end else begin
		if (soc_ethmac_writer_counter_ce) begin
			soc_ethmac_writer_counter <= (soc_ethmac_writer_counter + soc_ethmac_writer_increment);
		end
	end
	if (soc_ethmac_writer_slot_ce) begin
		soc_ethmac_writer_slot <= (soc_ethmac_writer_slot + 1'd1);
	end
	if (((soc_ethmac_writer_fifo_syncfifo_we & soc_ethmac_writer_fifo_syncfifo_writable) & (~soc_ethmac_writer_fifo_replace))) begin
		soc_ethmac_writer_fifo_produce <= (soc_ethmac_writer_fifo_produce + 1'd1);
	end
	if (soc_ethmac_writer_fifo_do_read) begin
		soc_ethmac_writer_fifo_consume <= (soc_ethmac_writer_fifo_consume + 1'd1);
	end
	if (((soc_ethmac_writer_fifo_syncfifo_we & soc_ethmac_writer_fifo_syncfifo_writable) & (~soc_ethmac_writer_fifo_replace))) begin
		if ((~soc_ethmac_writer_fifo_do_read)) begin
			soc_ethmac_writer_fifo_level <= (soc_ethmac_writer_fifo_level + 1'd1);
		end
	end else begin
		if (soc_ethmac_writer_fifo_do_read) begin
			soc_ethmac_writer_fifo_level <= (soc_ethmac_writer_fifo_level - 1'd1);
		end
	end
	vns_liteethmacsramwriter_state <= vns_liteethmacsramwriter_next_state;
	if (soc_ethmac_reader_counter_reset) begin
		soc_ethmac_reader_counter <= 1'd0;
	end else begin
		if (soc_ethmac_reader_counter_ce) begin
			soc_ethmac_reader_counter <= (soc_ethmac_reader_counter + 3'd4);
		end
	end
	if (soc_ethmac_reader_done_clear) begin
		soc_ethmac_reader_done_pending <= 1'd0;
	end
	if (soc_ethmac_reader_done_trigger) begin
		soc_ethmac_reader_done_pending <= 1'd1;
	end
	if (((soc_ethmac_reader_fifo_syncfifo_we & soc_ethmac_reader_fifo_syncfifo_writable) & (~soc_ethmac_reader_fifo_replace))) begin
		soc_ethmac_reader_fifo_produce <= (soc_ethmac_reader_fifo_produce + 1'd1);
	end
	if (soc_ethmac_reader_fifo_do_read) begin
		soc_ethmac_reader_fifo_consume <= (soc_ethmac_reader_fifo_consume + 1'd1);
	end
	if (((soc_ethmac_reader_fifo_syncfifo_we & soc_ethmac_reader_fifo_syncfifo_writable) & (~soc_ethmac_reader_fifo_replace))) begin
		if ((~soc_ethmac_reader_fifo_do_read)) begin
			soc_ethmac_reader_fifo_level <= (soc_ethmac_reader_fifo_level + 1'd1);
		end
	end else begin
		if (soc_ethmac_reader_fifo_do_read) begin
			soc_ethmac_reader_fifo_level <= (soc_ethmac_reader_fifo_level - 1'd1);
		end
	end
	vns_liteethmacsramreader_state <= vns_liteethmacsramreader_next_state;
	soc_ethmac_sram0_bus_ack0 <= 1'd0;
	if (((soc_ethmac_sram0_bus_cyc0 & soc_ethmac_sram0_bus_stb0) & (~soc_ethmac_sram0_bus_ack0))) begin
		soc_ethmac_sram0_bus_ack0 <= 1'd1;
	end
	soc_ethmac_sram1_bus_ack0 <= 1'd0;
	if (((soc_ethmac_sram1_bus_cyc0 & soc_ethmac_sram1_bus_stb0) & (~soc_ethmac_sram1_bus_ack0))) begin
		soc_ethmac_sram1_bus_ack0 <= 1'd1;
	end
	soc_ethmac_sram0_bus_ack1 <= 1'd0;
	if (((soc_ethmac_sram0_bus_cyc1 & soc_ethmac_sram0_bus_stb1) & (~soc_ethmac_sram0_bus_ack1))) begin
		soc_ethmac_sram0_bus_ack1 <= 1'd1;
	end
	soc_ethmac_sram1_bus_ack1 <= 1'd0;
	if (((soc_ethmac_sram1_bus_cyc1 & soc_ethmac_sram1_bus_stb1) & (~soc_ethmac_sram1_bus_ack1))) begin
		soc_ethmac_sram1_bus_ack1 <= 1'd1;
	end
	soc_ethmac_slave_sel_r <= soc_ethmac_slave_sel;
	soc_edid_sda_drv_reg <= soc_edid_sda_drv;
	{soc_edid_samp_carry, soc_edid_samp_count} <= (soc_edid_samp_count + 1'd1);
	if (soc_edid_samp_carry) begin
		soc_edid_scl_i <= soc_edid_scl_raw;
		soc_edid_sda_i <= soc_edid_sda_raw;
	end
	soc_edid_scl_r <= soc_edid_scl_i;
	soc_edid_sda_r <= soc_edid_sda_i;
	if (soc_edid_start) begin
		soc_edid_counter <= 1'd0;
	end
	if (soc_edid_scl_rising) begin
		if ((soc_edid_counter == 4'd8)) begin
			soc_edid_counter <= 1'd0;
		end else begin
			soc_edid_counter <= (soc_edid_counter + 1'd1);
			soc_edid_din <= {soc_edid_din[6:0], soc_edid_sda_i};
		end
	end
	if (soc_edid_update_is_read) begin
		soc_edid_is_read <= soc_edid_din[0];
	end
	if (soc_edid_oc_load) begin
		soc_edid_offset_counter <= soc_edid_din;
	end else begin
		if (soc_edid_oc_inc) begin
			soc_edid_offset_counter <= (soc_edid_offset_counter + 1'd1);
		end
	end
	if (soc_edid_data_drv_en) begin
		soc_edid_data_drv <= 1'd1;
	end else begin
		if (soc_edid_data_drv_stop) begin
			soc_edid_data_drv <= 1'd0;
		end
	end
	if (soc_edid_data_drv_en) begin
		case (soc_edid_counter)
			1'd0: begin
				soc_edid_data_bit <= soc_edid_dat_r[7];
			end
			1'd1: begin
				soc_edid_data_bit <= soc_edid_dat_r[6];
			end
			2'd2: begin
				soc_edid_data_bit <= soc_edid_dat_r[5];
			end
			2'd3: begin
				soc_edid_data_bit <= soc_edid_dat_r[4];
			end
			3'd4: begin
				soc_edid_data_bit <= soc_edid_dat_r[3];
			end
			3'd5: begin
				soc_edid_data_bit <= soc_edid_dat_r[2];
			end
			3'd6: begin
				soc_edid_data_bit <= soc_edid_dat_r[1];
			end
			default: begin
				soc_edid_data_bit <= soc_edid_dat_r[0];
			end
		endcase
	end
	vns_edid_state <= vns_edid_next_state;
	if ((soc_mmcm_read_re | soc_mmcm_write_re)) begin
		soc_mmcm_drdy_status <= 1'd0;
	end else begin
		if (soc_mmcm_drdy) begin
			soc_mmcm_drdy_status <= 1'd1;
		end
	end
	if (soc_s7datacapture0_do_delay_rst_i) begin
		soc_s7datacapture0_do_delay_rst_toggle_i <= (~soc_s7datacapture0_do_delay_rst_toggle_i);
	end
	if (soc_s7datacapture0_do_delay_master_inc_i) begin
		soc_s7datacapture0_do_delay_master_inc_toggle_i <= (~soc_s7datacapture0_do_delay_master_inc_toggle_i);
	end
	if (soc_s7datacapture0_do_delay_master_dec_i) begin
		soc_s7datacapture0_do_delay_master_dec_toggle_i <= (~soc_s7datacapture0_do_delay_master_dec_toggle_i);
	end
	if (soc_s7datacapture0_do_delay_slave_inc_i) begin
		soc_s7datacapture0_do_delay_slave_inc_toggle_i <= (~soc_s7datacapture0_do_delay_slave_inc_toggle_i);
	end
	if (soc_s7datacapture0_do_delay_slave_dec_i) begin
		soc_s7datacapture0_do_delay_slave_dec_toggle_i <= (~soc_s7datacapture0_do_delay_slave_dec_toggle_i);
	end
	if (soc_s7datacapture0_do_reset_lateness_i) begin
		soc_s7datacapture0_do_reset_lateness_toggle_i <= (~soc_s7datacapture0_do_reset_lateness_toggle_i);
	end
	if (soc_wer0_o) begin
		soc_wer0_wer_counter_sys <= soc_wer0_wer_counter_r;
	end
	if (soc_wer0_update_re) begin
		soc_wer0_status <= soc_wer0_wer_counter_sys;
	end
	soc_wer0_toggle_o_r <= soc_wer0_toggle_o;
	if (soc_s7datacapture1_do_delay_rst_i) begin
		soc_s7datacapture1_do_delay_rst_toggle_i <= (~soc_s7datacapture1_do_delay_rst_toggle_i);
	end
	if (soc_s7datacapture1_do_delay_master_inc_i) begin
		soc_s7datacapture1_do_delay_master_inc_toggle_i <= (~soc_s7datacapture1_do_delay_master_inc_toggle_i);
	end
	if (soc_s7datacapture1_do_delay_master_dec_i) begin
		soc_s7datacapture1_do_delay_master_dec_toggle_i <= (~soc_s7datacapture1_do_delay_master_dec_toggle_i);
	end
	if (soc_s7datacapture1_do_delay_slave_inc_i) begin
		soc_s7datacapture1_do_delay_slave_inc_toggle_i <= (~soc_s7datacapture1_do_delay_slave_inc_toggle_i);
	end
	if (soc_s7datacapture1_do_delay_slave_dec_i) begin
		soc_s7datacapture1_do_delay_slave_dec_toggle_i <= (~soc_s7datacapture1_do_delay_slave_dec_toggle_i);
	end
	if (soc_s7datacapture1_do_reset_lateness_i) begin
		soc_s7datacapture1_do_reset_lateness_toggle_i <= (~soc_s7datacapture1_do_reset_lateness_toggle_i);
	end
	if (soc_wer1_o) begin
		soc_wer1_wer_counter_sys <= soc_wer1_wer_counter_r;
	end
	if (soc_wer1_update_re) begin
		soc_wer1_status <= soc_wer1_wer_counter_sys;
	end
	soc_wer1_toggle_o_r <= soc_wer1_toggle_o;
	if (soc_s7datacapture2_do_delay_rst_i) begin
		soc_s7datacapture2_do_delay_rst_toggle_i <= (~soc_s7datacapture2_do_delay_rst_toggle_i);
	end
	if (soc_s7datacapture2_do_delay_master_inc_i) begin
		soc_s7datacapture2_do_delay_master_inc_toggle_i <= (~soc_s7datacapture2_do_delay_master_inc_toggle_i);
	end
	if (soc_s7datacapture2_do_delay_master_dec_i) begin
		soc_s7datacapture2_do_delay_master_dec_toggle_i <= (~soc_s7datacapture2_do_delay_master_dec_toggle_i);
	end
	if (soc_s7datacapture2_do_delay_slave_inc_i) begin
		soc_s7datacapture2_do_delay_slave_inc_toggle_i <= (~soc_s7datacapture2_do_delay_slave_inc_toggle_i);
	end
	if (soc_s7datacapture2_do_delay_slave_dec_i) begin
		soc_s7datacapture2_do_delay_slave_dec_toggle_i <= (~soc_s7datacapture2_do_delay_slave_dec_toggle_i);
	end
	if (soc_s7datacapture2_do_reset_lateness_i) begin
		soc_s7datacapture2_do_reset_lateness_toggle_i <= (~soc_s7datacapture2_do_reset_lateness_toggle_i);
	end
	if (soc_wer2_o) begin
		soc_wer2_wer_counter_sys <= soc_wer2_wer_counter_r;
	end
	if (soc_wer2_update_re) begin
		soc_wer2_status <= soc_wer2_wer_counter_sys;
	end
	soc_wer2_toggle_o_r <= soc_wer2_toggle_o;
	if (soc_frame_overflow_re) begin
		soc_frame_overflow_mask <= 1'd1;
	end else begin
		if (soc_frame_overflow_reset_ack_o) begin
			soc_frame_overflow_mask <= 1'd0;
		end
	end
	soc_frame_fifo_graycounter1_q_binary <= soc_frame_fifo_graycounter1_q_next_binary;
	soc_frame_fifo_graycounter1_q <= soc_frame_fifo_graycounter1_q_next;
	if (soc_frame_overflow_reset_i) begin
		soc_frame_overflow_reset_toggle_i <= (~soc_frame_overflow_reset_toggle_i);
	end
	soc_frame_overflow_reset_ack_toggle_o_r <= soc_frame_overflow_reset_ack_toggle_o;
	if (soc_dma_reset_words) begin
		soc_dma_current_address <= soc_dma_slot_array_address;
		soc_dma_mwords_remaining <= soc_dma_frame_size_storage;
	end else begin
		if (soc_dma_count_word) begin
			soc_dma_current_address <= (soc_dma_current_address + 1'd1);
			soc_dma_mwords_remaining <= (soc_dma_mwords_remaining - 1'd1);
		end
	end
	if (soc_dma_slot_array_change_slot) begin
		if (soc_dma_slot_array_slot1_address_valid) begin
			soc_dma_slot_array_current_slot <= 1'd1;
		end
		if (soc_dma_slot_array_slot0_address_valid) begin
			soc_dma_slot_array_current_slot <= 1'd0;
		end
	end
	if (((soc_dma_fifo_syncfifo_we & soc_dma_fifo_syncfifo_writable) & (~soc_dma_fifo_replace))) begin
		soc_dma_fifo_produce <= (soc_dma_fifo_produce + 1'd1);
	end
	if (soc_dma_fifo_do_read) begin
		soc_dma_fifo_consume <= (soc_dma_fifo_consume + 1'd1);
	end
	if (((soc_dma_fifo_syncfifo_we & soc_dma_fifo_syncfifo_writable) & (~soc_dma_fifo_replace))) begin
		if ((~soc_dma_fifo_do_read)) begin
			soc_dma_fifo_level <= (soc_dma_fifo_level + 1'd1);
		end
	end else begin
		if (soc_dma_fifo_do_read) begin
			soc_dma_fifo_level <= (soc_dma_fifo_level - 1'd1);
		end
	end
	vns_dma_state <= vns_dma_next_state;
	if (soc_hdmi_in0_freq_period_done) begin
		soc_hdmi_in0_freq_period_counter <= 1'd0;
	end else begin
		soc_hdmi_in0_freq_period_counter <= (soc_hdmi_in0_freq_period_counter + 1'd1);
	end
	soc_hdmi_in0_freq_gray_decoder_o <= soc_hdmi_in0_freq_gray_decoder_o_comb;
	soc_hdmi_in0_freq_sampler_i_d <= soc_hdmi_in0_freq_sampler_i;
	if (soc_hdmi_in0_freq_sampler_latch) begin
		soc_hdmi_in0_freq_sampler_counter <= 1'd0;
		soc_hdmi_in0_freq_sampler_o <= soc_hdmi_in0_freq_sampler_counter;
	end else begin
		soc_hdmi_in0_freq_sampler_counter <= (soc_hdmi_in0_freq_sampler_counter + soc_hdmi_in0_freq_sampler_inc);
	end
	soc_hdmi_out0_core_initiator_cdc_graycounter0_q_binary <= soc_hdmi_out0_core_initiator_cdc_graycounter0_q_next_binary;
	soc_hdmi_out0_core_initiator_cdc_graycounter0_q <= soc_hdmi_out0_core_initiator_cdc_graycounter0_q_next;
	if (soc_hdmi_out0_core_i) begin
		soc_hdmi_out0_core_toggle_i <= (~soc_hdmi_out0_core_toggle_i);
	end
	if ((soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_read_re | soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_write_re)) begin
		soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy_status <= 1'd0;
	end else begin
		if (soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy) begin
			soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy_status <= 1'd1;
		end
	end
	case (vns_videosoc_grant)
		1'd0: begin
			if ((~vns_videosoc_request[0])) begin
				if (vns_videosoc_request[1]) begin
					vns_videosoc_grant <= 1'd1;
				end else begin
					if (vns_videosoc_request[2]) begin
						vns_videosoc_grant <= 2'd2;
					end
				end
			end
		end
		1'd1: begin
			if ((~vns_videosoc_request[1])) begin
				if (vns_videosoc_request[2]) begin
					vns_videosoc_grant <= 2'd2;
				end else begin
					if (vns_videosoc_request[0]) begin
						vns_videosoc_grant <= 1'd0;
					end
				end
			end
		end
		2'd2: begin
			if ((~vns_videosoc_request[2])) begin
				if (vns_videosoc_request[0]) begin
					vns_videosoc_grant <= 1'd0;
				end else begin
					if (vns_videosoc_request[1]) begin
						vns_videosoc_grant <= 1'd1;
					end
				end
			end
		end
	endcase
	vns_videosoc_slave_sel_r <= vns_videosoc_slave_sel;
	vns_videosoc_interface0_bank_bus_dat_r <= 1'd0;
	if (vns_videosoc_csrbank0_sel) begin
		case (vns_videosoc_interface0_bank_bus_adr[1:0])
			1'd0: begin
				vns_videosoc_interface0_bank_bus_dat_r <= vns_videosoc_csrbank0_dly_sel0_w;
			end
			1'd1: begin
				vns_videosoc_interface0_bank_bus_dat_r <= soc_videosoc_ddrphy_rdly_dq_rst_w;
			end
			2'd2: begin
				vns_videosoc_interface0_bank_bus_dat_r <= soc_videosoc_ddrphy_rdly_dq_inc_w;
			end
			2'd3: begin
				vns_videosoc_interface0_bank_bus_dat_r <= soc_videosoc_ddrphy_rdly_dq_bitslip_w;
			end
		endcase
	end
	if (vns_videosoc_csrbank0_dly_sel0_re) begin
		soc_videosoc_ddrphy_storage_full[1:0] <= vns_videosoc_csrbank0_dly_sel0_r;
	end
	soc_videosoc_ddrphy_re <= vns_videosoc_csrbank0_dly_sel0_re;
	vns_videosoc_interface1_bank_bus_dat_r <= 1'd0;
	if (vns_videosoc_csrbank1_sel) begin
		case (vns_videosoc_interface1_bank_bus_adr[4:0])
			1'd0: begin
				vns_videosoc_interface1_bank_bus_dat_r <= vns_videosoc_csrbank1_sram_writer_slot_w;
			end
			1'd1: begin
				vns_videosoc_interface1_bank_bus_dat_r <= vns_videosoc_csrbank1_sram_writer_length3_w;
			end
			2'd2: begin
				vns_videosoc_interface1_bank_bus_dat_r <= vns_videosoc_csrbank1_sram_writer_length2_w;
			end
			2'd3: begin
				vns_videosoc_interface1_bank_bus_dat_r <= vns_videosoc_csrbank1_sram_writer_length1_w;
			end
			3'd4: begin
				vns_videosoc_interface1_bank_bus_dat_r <= vns_videosoc_csrbank1_sram_writer_length0_w;
			end
			3'd5: begin
				vns_videosoc_interface1_bank_bus_dat_r <= soc_ethmac_writer_status_w;
			end
			3'd6: begin
				vns_videosoc_interface1_bank_bus_dat_r <= soc_ethmac_writer_pending_w;
			end
			3'd7: begin
				vns_videosoc_interface1_bank_bus_dat_r <= vns_videosoc_csrbank1_sram_writer_ev_enable0_w;
			end
			4'd8: begin
				vns_videosoc_interface1_bank_bus_dat_r <= soc_ethmac_reader_start_w;
			end
			4'd9: begin
				vns_videosoc_interface1_bank_bus_dat_r <= vns_videosoc_csrbank1_sram_reader_ready_w;
			end
			4'd10: begin
				vns_videosoc_interface1_bank_bus_dat_r <= vns_videosoc_csrbank1_sram_reader_slot0_w;
			end
			4'd11: begin
				vns_videosoc_interface1_bank_bus_dat_r <= vns_videosoc_csrbank1_sram_reader_length1_w;
			end
			4'd12: begin
				vns_videosoc_interface1_bank_bus_dat_r <= vns_videosoc_csrbank1_sram_reader_length0_w;
			end
			4'd13: begin
				vns_videosoc_interface1_bank_bus_dat_r <= soc_ethmac_reader_eventmanager_status_w;
			end
			4'd14: begin
				vns_videosoc_interface1_bank_bus_dat_r <= soc_ethmac_reader_eventmanager_pending_w;
			end
			4'd15: begin
				vns_videosoc_interface1_bank_bus_dat_r <= vns_videosoc_csrbank1_sram_reader_ev_enable0_w;
			end
			5'd16: begin
				vns_videosoc_interface1_bank_bus_dat_r <= vns_videosoc_csrbank1_preamble_crc_w;
			end
		endcase
	end
	if (vns_videosoc_csrbank1_sram_writer_ev_enable0_re) begin
		soc_ethmac_writer_storage_full <= vns_videosoc_csrbank1_sram_writer_ev_enable0_r;
	end
	soc_ethmac_writer_re <= vns_videosoc_csrbank1_sram_writer_ev_enable0_re;
	if (vns_videosoc_csrbank1_sram_reader_slot0_re) begin
		soc_ethmac_reader_slot_storage_full <= vns_videosoc_csrbank1_sram_reader_slot0_r;
	end
	soc_ethmac_reader_slot_re <= vns_videosoc_csrbank1_sram_reader_slot0_re;
	if (vns_videosoc_csrbank1_sram_reader_length1_re) begin
		soc_ethmac_reader_length_storage_full[10:8] <= vns_videosoc_csrbank1_sram_reader_length1_r;
	end
	if (vns_videosoc_csrbank1_sram_reader_length0_re) begin
		soc_ethmac_reader_length_storage_full[7:0] <= vns_videosoc_csrbank1_sram_reader_length0_r;
	end
	soc_ethmac_reader_length_re <= vns_videosoc_csrbank1_sram_reader_length0_re;
	if (vns_videosoc_csrbank1_sram_reader_ev_enable0_re) begin
		soc_ethmac_reader_eventmanager_storage_full <= vns_videosoc_csrbank1_sram_reader_ev_enable0_r;
	end
	soc_ethmac_reader_eventmanager_re <= vns_videosoc_csrbank1_sram_reader_ev_enable0_re;
	vns_videosoc_interface2_bank_bus_dat_r <= 1'd0;
	if (vns_videosoc_csrbank2_sel) begin
		case (vns_videosoc_interface2_bank_bus_adr[1:0])
			1'd0: begin
				vns_videosoc_interface2_bank_bus_dat_r <= vns_videosoc_csrbank2_crg_reset0_w;
			end
			1'd1: begin
				vns_videosoc_interface2_bank_bus_dat_r <= vns_videosoc_csrbank2_mdio_w0_w;
			end
			2'd2: begin
				vns_videosoc_interface2_bank_bus_dat_r <= vns_videosoc_csrbank2_mdio_r_w;
			end
		endcase
	end
	if (vns_videosoc_csrbank2_crg_reset0_re) begin
		soc_ethphy_reset_storage_full <= vns_videosoc_csrbank2_crg_reset0_r;
	end
	soc_ethphy_reset_re <= vns_videosoc_csrbank2_crg_reset0_re;
	if (vns_videosoc_csrbank2_mdio_w0_re) begin
		soc_ethphy_storage_full[2:0] <= vns_videosoc_csrbank2_mdio_w0_r;
	end
	soc_ethphy_re <= vns_videosoc_csrbank2_mdio_w0_re;
	vns_videosoc_sel_r <= vns_videosoc_sel;
	vns_videosoc_interface3_bank_bus_dat_r <= 1'd0;
	if (vns_videosoc_csrbank3_sel) begin
		case (vns_videosoc_interface3_bank_bus_adr[5:0])
			1'd0: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_edid_hpd_notif_w;
			end
			1'd1: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_edid_hpd_en0_w;
			end
			2'd2: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_clocking_mmcm_reset0_w;
			end
			2'd3: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_clocking_locked_w;
			end
			3'd4: begin
				vns_videosoc_interface3_bank_bus_dat_r <= soc_mmcm_read_w;
			end
			3'd5: begin
				vns_videosoc_interface3_bank_bus_dat_r <= soc_mmcm_write_w;
			end
			3'd6: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_clocking_mmcm_drdy_w;
			end
			3'd7: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_clocking_mmcm_adr0_w;
			end
			4'd8: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_clocking_mmcm_dat_w1_w;
			end
			4'd9: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_clocking_mmcm_dat_w0_w;
			end
			4'd10: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_clocking_mmcm_dat_r1_w;
			end
			4'd11: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_clocking_mmcm_dat_r0_w;
			end
			4'd12: begin
				vns_videosoc_interface3_bank_bus_dat_r <= soc_s7datacapture0_dly_ctl_w;
			end
			4'd13: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data0_cap_phase_w;
			end
			4'd14: begin
				vns_videosoc_interface3_bank_bus_dat_r <= soc_s7datacapture0_phase_reset_w;
			end
			4'd15: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data0_charsync_char_synced_w;
			end
			5'd16: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data0_charsync_ctl_pos_w;
			end
			5'd17: begin
				vns_videosoc_interface3_bank_bus_dat_r <= soc_wer0_update_w;
			end
			5'd18: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data0_wer_value2_w;
			end
			5'd19: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data0_wer_value1_w;
			end
			5'd20: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data0_wer_value0_w;
			end
			5'd21: begin
				vns_videosoc_interface3_bank_bus_dat_r <= soc_s7datacapture1_dly_ctl_w;
			end
			5'd22: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data1_cap_phase_w;
			end
			5'd23: begin
				vns_videosoc_interface3_bank_bus_dat_r <= soc_s7datacapture1_phase_reset_w;
			end
			5'd24: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data1_charsync_char_synced_w;
			end
			5'd25: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data1_charsync_ctl_pos_w;
			end
			5'd26: begin
				vns_videosoc_interface3_bank_bus_dat_r <= soc_wer1_update_w;
			end
			5'd27: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data1_wer_value2_w;
			end
			5'd28: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data1_wer_value1_w;
			end
			5'd29: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data1_wer_value0_w;
			end
			5'd30: begin
				vns_videosoc_interface3_bank_bus_dat_r <= soc_s7datacapture2_dly_ctl_w;
			end
			5'd31: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data2_cap_phase_w;
			end
			6'd32: begin
				vns_videosoc_interface3_bank_bus_dat_r <= soc_s7datacapture2_phase_reset_w;
			end
			6'd33: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data2_charsync_char_synced_w;
			end
			6'd34: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data2_charsync_ctl_pos_w;
			end
			6'd35: begin
				vns_videosoc_interface3_bank_bus_dat_r <= soc_wer2_update_w;
			end
			6'd36: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data2_wer_value2_w;
			end
			6'd37: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data2_wer_value1_w;
			end
			6'd38: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_data2_wer_value0_w;
			end
			6'd39: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_chansync_channels_synced_w;
			end
			6'd40: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_resdetection_hres1_w;
			end
			6'd41: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_resdetection_hres0_w;
			end
			6'd42: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_resdetection_vres1_w;
			end
			6'd43: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_resdetection_vres0_w;
			end
			6'd44: begin
				vns_videosoc_interface3_bank_bus_dat_r <= soc_frame_overflow_w;
			end
			6'd45: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_dma_frame_size3_w;
			end
			6'd46: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_dma_frame_size2_w;
			end
			6'd47: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_dma_frame_size1_w;
			end
			6'd48: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_dma_frame_size0_w;
			end
			6'd49: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_dma_slot0_status0_w;
			end
			6'd50: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_dma_slot0_address3_w;
			end
			6'd51: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_dma_slot0_address2_w;
			end
			6'd52: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_dma_slot0_address1_w;
			end
			6'd53: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_dma_slot0_address0_w;
			end
			6'd54: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_dma_slot1_status0_w;
			end
			6'd55: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_dma_slot1_address3_w;
			end
			6'd56: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_dma_slot1_address2_w;
			end
			6'd57: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_dma_slot1_address1_w;
			end
			6'd58: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_dma_slot1_address0_w;
			end
			6'd59: begin
				vns_videosoc_interface3_bank_bus_dat_r <= soc_dma_slot_array_status_w;
			end
			6'd60: begin
				vns_videosoc_interface3_bank_bus_dat_r <= soc_dma_slot_array_pending_w;
			end
			6'd61: begin
				vns_videosoc_interface3_bank_bus_dat_r <= vns_videosoc_csrbank3_dma_ev_enable0_w;
			end
		endcase
	end
	if (vns_videosoc_csrbank3_edid_hpd_en0_re) begin
		soc_edid_storage_full <= vns_videosoc_csrbank3_edid_hpd_en0_r;
	end
	soc_edid_re <= vns_videosoc_csrbank3_edid_hpd_en0_re;
	if (vns_videosoc_csrbank3_clocking_mmcm_reset0_re) begin
		soc_mmcm_reset_storage_full <= vns_videosoc_csrbank3_clocking_mmcm_reset0_r;
	end
	soc_mmcm_reset_re <= vns_videosoc_csrbank3_clocking_mmcm_reset0_re;
	if (vns_videosoc_csrbank3_clocking_mmcm_adr0_re) begin
		soc_mmcm_adr_storage_full[6:0] <= vns_videosoc_csrbank3_clocking_mmcm_adr0_r;
	end
	soc_mmcm_adr_re <= vns_videosoc_csrbank3_clocking_mmcm_adr0_re;
	if (vns_videosoc_csrbank3_clocking_mmcm_dat_w1_re) begin
		soc_mmcm_dat_w_storage_full[15:8] <= vns_videosoc_csrbank3_clocking_mmcm_dat_w1_r;
	end
	if (vns_videosoc_csrbank3_clocking_mmcm_dat_w0_re) begin
		soc_mmcm_dat_w_storage_full[7:0] <= vns_videosoc_csrbank3_clocking_mmcm_dat_w0_r;
	end
	soc_mmcm_dat_w_re <= vns_videosoc_csrbank3_clocking_mmcm_dat_w0_re;
	if (vns_videosoc_csrbank3_dma_frame_size3_re) begin
		soc_dma_frame_size_storage_full[28:24] <= vns_videosoc_csrbank3_dma_frame_size3_r;
	end
	if (vns_videosoc_csrbank3_dma_frame_size2_re) begin
		soc_dma_frame_size_storage_full[23:16] <= vns_videosoc_csrbank3_dma_frame_size2_r;
	end
	if (vns_videosoc_csrbank3_dma_frame_size1_re) begin
		soc_dma_frame_size_storage_full[15:8] <= vns_videosoc_csrbank3_dma_frame_size1_r;
	end
	if (vns_videosoc_csrbank3_dma_frame_size0_re) begin
		soc_dma_frame_size_storage_full[7:0] <= vns_videosoc_csrbank3_dma_frame_size0_r;
	end
	soc_dma_frame_size_re <= vns_videosoc_csrbank3_dma_frame_size0_re;
	if (soc_dma_slot_array_slot0_status_we) begin
		soc_dma_slot_array_slot0_status_storage_full <= (soc_dma_slot_array_slot0_status_dat_w <<< 1'd0);
	end
	if (vns_videosoc_csrbank3_dma_slot0_status0_re) begin
		soc_dma_slot_array_slot0_status_storage_full[1:0] <= vns_videosoc_csrbank3_dma_slot0_status0_r;
	end
	soc_dma_slot_array_slot0_status_re <= vns_videosoc_csrbank3_dma_slot0_status0_re;
	if (soc_dma_slot_array_slot0_address_we) begin
		soc_dma_slot_array_slot0_address_storage_full <= (soc_dma_slot_array_slot0_address_dat_w <<< 3'd4);
	end
	if (vns_videosoc_csrbank3_dma_slot0_address3_re) begin
		soc_dma_slot_array_slot0_address_storage_full[28:24] <= vns_videosoc_csrbank3_dma_slot0_address3_r;
	end
	if (vns_videosoc_csrbank3_dma_slot0_address2_re) begin
		soc_dma_slot_array_slot0_address_storage_full[23:16] <= vns_videosoc_csrbank3_dma_slot0_address2_r;
	end
	if (vns_videosoc_csrbank3_dma_slot0_address1_re) begin
		soc_dma_slot_array_slot0_address_storage_full[15:8] <= vns_videosoc_csrbank3_dma_slot0_address1_r;
	end
	if (vns_videosoc_csrbank3_dma_slot0_address0_re) begin
		soc_dma_slot_array_slot0_address_storage_full[7:0] <= vns_videosoc_csrbank3_dma_slot0_address0_r;
	end
	soc_dma_slot_array_slot0_address_re <= vns_videosoc_csrbank3_dma_slot0_address0_re;
	if (soc_dma_slot_array_slot1_status_we) begin
		soc_dma_slot_array_slot1_status_storage_full <= (soc_dma_slot_array_slot1_status_dat_w <<< 1'd0);
	end
	if (vns_videosoc_csrbank3_dma_slot1_status0_re) begin
		soc_dma_slot_array_slot1_status_storage_full[1:0] <= vns_videosoc_csrbank3_dma_slot1_status0_r;
	end
	soc_dma_slot_array_slot1_status_re <= vns_videosoc_csrbank3_dma_slot1_status0_re;
	if (soc_dma_slot_array_slot1_address_we) begin
		soc_dma_slot_array_slot1_address_storage_full <= (soc_dma_slot_array_slot1_address_dat_w <<< 3'd4);
	end
	if (vns_videosoc_csrbank3_dma_slot1_address3_re) begin
		soc_dma_slot_array_slot1_address_storage_full[28:24] <= vns_videosoc_csrbank3_dma_slot1_address3_r;
	end
	if (vns_videosoc_csrbank3_dma_slot1_address2_re) begin
		soc_dma_slot_array_slot1_address_storage_full[23:16] <= vns_videosoc_csrbank3_dma_slot1_address2_r;
	end
	if (vns_videosoc_csrbank3_dma_slot1_address1_re) begin
		soc_dma_slot_array_slot1_address_storage_full[15:8] <= vns_videosoc_csrbank3_dma_slot1_address1_r;
	end
	if (vns_videosoc_csrbank3_dma_slot1_address0_re) begin
		soc_dma_slot_array_slot1_address_storage_full[7:0] <= vns_videosoc_csrbank3_dma_slot1_address0_r;
	end
	soc_dma_slot_array_slot1_address_re <= vns_videosoc_csrbank3_dma_slot1_address0_re;
	if (vns_videosoc_csrbank3_dma_ev_enable0_re) begin
		soc_dma_slot_array_storage_full[1:0] <= vns_videosoc_csrbank3_dma_ev_enable0_r;
	end
	soc_dma_slot_array_re <= vns_videosoc_csrbank3_dma_ev_enable0_re;
	vns_videosoc_interface4_bank_bus_dat_r <= 1'd0;
	if (vns_videosoc_csrbank4_sel) begin
		case (vns_videosoc_interface4_bank_bus_adr[1:0])
			1'd0: begin
				vns_videosoc_interface4_bank_bus_dat_r <= vns_videosoc_csrbank4_value3_w;
			end
			1'd1: begin
				vns_videosoc_interface4_bank_bus_dat_r <= vns_videosoc_csrbank4_value2_w;
			end
			2'd2: begin
				vns_videosoc_interface4_bank_bus_dat_r <= vns_videosoc_csrbank4_value1_w;
			end
			2'd3: begin
				vns_videosoc_interface4_bank_bus_dat_r <= vns_videosoc_csrbank4_value0_w;
			end
		endcase
	end
	vns_videosoc_interface5_bank_bus_dat_r <= 1'd0;
	if (vns_videosoc_csrbank5_sel) begin
		case (vns_videosoc_interface5_bank_bus_adr[5:0])
			1'd0: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_underflow_enable0_w;
			end
			1'd1: begin
				vns_videosoc_interface5_bank_bus_dat_r <= soc_hdmi_out0_core_underflow_update_underflow_update_w;
			end
			2'd2: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_underflow_counter3_w;
			end
			2'd3: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_underflow_counter2_w;
			end
			3'd4: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_underflow_counter1_w;
			end
			3'd5: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_underflow_counter0_w;
			end
			3'd6: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_enable0_w;
			end
			3'd7: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_hres1_w;
			end
			4'd8: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_hres0_w;
			end
			4'd9: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_hsync_start1_w;
			end
			4'd10: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_hsync_start0_w;
			end
			4'd11: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_hsync_end1_w;
			end
			4'd12: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_hsync_end0_w;
			end
			4'd13: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_hscan1_w;
			end
			4'd14: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_hscan0_w;
			end
			4'd15: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_vres1_w;
			end
			5'd16: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_vres0_w;
			end
			5'd17: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_vsync_start1_w;
			end
			5'd18: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_vsync_start0_w;
			end
			5'd19: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_vsync_end1_w;
			end
			5'd20: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_vsync_end0_w;
			end
			5'd21: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_vscan1_w;
			end
			5'd22: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_vscan0_w;
			end
			5'd23: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_base3_w;
			end
			5'd24: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_base2_w;
			end
			5'd25: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_base1_w;
			end
			5'd26: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_base0_w;
			end
			5'd27: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_length3_w;
			end
			5'd28: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_length2_w;
			end
			5'd29: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_length1_w;
			end
			5'd30: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_core_initiator_length0_w;
			end
			5'd31: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_driver_clocking_mmcm_reset0_w;
			end
			6'd32: begin
				vns_videosoc_interface5_bank_bus_dat_r <= soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_read_w;
			end
			6'd33: begin
				vns_videosoc_interface5_bank_bus_dat_r <= soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_write_w;
			end
			6'd34: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_driver_clocking_mmcm_drdy_w;
			end
			6'd35: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_driver_clocking_mmcm_adr0_w;
			end
			6'd36: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w1_w;
			end
			6'd37: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w0_w;
			end
			6'd38: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_driver_clocking_mmcm_dat_r1_w;
			end
			6'd39: begin
				vns_videosoc_interface5_bank_bus_dat_r <= vns_videosoc_csrbank5_driver_clocking_mmcm_dat_r0_w;
			end
		endcase
	end
	if (vns_videosoc_csrbank5_core_underflow_enable0_re) begin
		soc_hdmi_out0_core_underflow_enable_storage_full <= vns_videosoc_csrbank5_core_underflow_enable0_r;
	end
	soc_hdmi_out0_core_underflow_enable_re <= vns_videosoc_csrbank5_core_underflow_enable0_re;
	if (vns_videosoc_csrbank5_core_initiator_enable0_re) begin
		soc_hdmi_out0_core_initiator_enable_storage_full <= vns_videosoc_csrbank5_core_initiator_enable0_r;
	end
	soc_hdmi_out0_core_initiator_enable_re <= vns_videosoc_csrbank5_core_initiator_enable0_re;
	if (vns_videosoc_csrbank5_core_initiator_hres1_re) begin
		vns_videosoc_csrbank5_core_initiator_hres_backstore[3:0] <= vns_videosoc_csrbank5_core_initiator_hres1_r;
	end
	if (vns_videosoc_csrbank5_core_initiator_hres0_re) begin
		soc_hdmi_out0_core_initiator_csrstorage0_storage_full <= {vns_videosoc_csrbank5_core_initiator_hres_backstore, vns_videosoc_csrbank5_core_initiator_hres0_r};
	end
	soc_hdmi_out0_core_initiator_csrstorage0_re <= vns_videosoc_csrbank5_core_initiator_hres0_re;
	if (vns_videosoc_csrbank5_core_initiator_hsync_start1_re) begin
		vns_videosoc_csrbank5_core_initiator_hsync_start_backstore[3:0] <= vns_videosoc_csrbank5_core_initiator_hsync_start1_r;
	end
	if (vns_videosoc_csrbank5_core_initiator_hsync_start0_re) begin
		soc_hdmi_out0_core_initiator_csrstorage1_storage_full <= {vns_videosoc_csrbank5_core_initiator_hsync_start_backstore, vns_videosoc_csrbank5_core_initiator_hsync_start0_r};
	end
	soc_hdmi_out0_core_initiator_csrstorage1_re <= vns_videosoc_csrbank5_core_initiator_hsync_start0_re;
	if (vns_videosoc_csrbank5_core_initiator_hsync_end1_re) begin
		vns_videosoc_csrbank5_core_initiator_hsync_end_backstore[3:0] <= vns_videosoc_csrbank5_core_initiator_hsync_end1_r;
	end
	if (vns_videosoc_csrbank5_core_initiator_hsync_end0_re) begin
		soc_hdmi_out0_core_initiator_csrstorage2_storage_full <= {vns_videosoc_csrbank5_core_initiator_hsync_end_backstore, vns_videosoc_csrbank5_core_initiator_hsync_end0_r};
	end
	soc_hdmi_out0_core_initiator_csrstorage2_re <= vns_videosoc_csrbank5_core_initiator_hsync_end0_re;
	if (vns_videosoc_csrbank5_core_initiator_hscan1_re) begin
		vns_videosoc_csrbank5_core_initiator_hscan_backstore[3:0] <= vns_videosoc_csrbank5_core_initiator_hscan1_r;
	end
	if (vns_videosoc_csrbank5_core_initiator_hscan0_re) begin
		soc_hdmi_out0_core_initiator_csrstorage3_storage_full <= {vns_videosoc_csrbank5_core_initiator_hscan_backstore, vns_videosoc_csrbank5_core_initiator_hscan0_r};
	end
	soc_hdmi_out0_core_initiator_csrstorage3_re <= vns_videosoc_csrbank5_core_initiator_hscan0_re;
	if (vns_videosoc_csrbank5_core_initiator_vres1_re) begin
		vns_videosoc_csrbank5_core_initiator_vres_backstore[3:0] <= vns_videosoc_csrbank5_core_initiator_vres1_r;
	end
	if (vns_videosoc_csrbank5_core_initiator_vres0_re) begin
		soc_hdmi_out0_core_initiator_csrstorage4_storage_full <= {vns_videosoc_csrbank5_core_initiator_vres_backstore, vns_videosoc_csrbank5_core_initiator_vres0_r};
	end
	soc_hdmi_out0_core_initiator_csrstorage4_re <= vns_videosoc_csrbank5_core_initiator_vres0_re;
	if (vns_videosoc_csrbank5_core_initiator_vsync_start1_re) begin
		vns_videosoc_csrbank5_core_initiator_vsync_start_backstore[3:0] <= vns_videosoc_csrbank5_core_initiator_vsync_start1_r;
	end
	if (vns_videosoc_csrbank5_core_initiator_vsync_start0_re) begin
		soc_hdmi_out0_core_initiator_csrstorage5_storage_full <= {vns_videosoc_csrbank5_core_initiator_vsync_start_backstore, vns_videosoc_csrbank5_core_initiator_vsync_start0_r};
	end
	soc_hdmi_out0_core_initiator_csrstorage5_re <= vns_videosoc_csrbank5_core_initiator_vsync_start0_re;
	if (vns_videosoc_csrbank5_core_initiator_vsync_end1_re) begin
		vns_videosoc_csrbank5_core_initiator_vsync_end_backstore[3:0] <= vns_videosoc_csrbank5_core_initiator_vsync_end1_r;
	end
	if (vns_videosoc_csrbank5_core_initiator_vsync_end0_re) begin
		soc_hdmi_out0_core_initiator_csrstorage6_storage_full <= {vns_videosoc_csrbank5_core_initiator_vsync_end_backstore, vns_videosoc_csrbank5_core_initiator_vsync_end0_r};
	end
	soc_hdmi_out0_core_initiator_csrstorage6_re <= vns_videosoc_csrbank5_core_initiator_vsync_end0_re;
	if (vns_videosoc_csrbank5_core_initiator_vscan1_re) begin
		vns_videosoc_csrbank5_core_initiator_vscan_backstore[3:0] <= vns_videosoc_csrbank5_core_initiator_vscan1_r;
	end
	if (vns_videosoc_csrbank5_core_initiator_vscan0_re) begin
		soc_hdmi_out0_core_initiator_csrstorage7_storage_full <= {vns_videosoc_csrbank5_core_initiator_vscan_backstore, vns_videosoc_csrbank5_core_initiator_vscan0_r};
	end
	soc_hdmi_out0_core_initiator_csrstorage7_re <= vns_videosoc_csrbank5_core_initiator_vscan0_re;
	if (vns_videosoc_csrbank5_core_initiator_base3_re) begin
		vns_videosoc_csrbank5_core_initiator_base_backstore[23:16] <= vns_videosoc_csrbank5_core_initiator_base3_r;
	end
	if (vns_videosoc_csrbank5_core_initiator_base2_re) begin
		vns_videosoc_csrbank5_core_initiator_base_backstore[15:8] <= vns_videosoc_csrbank5_core_initiator_base2_r;
	end
	if (vns_videosoc_csrbank5_core_initiator_base1_re) begin
		vns_videosoc_csrbank5_core_initiator_base_backstore[7:0] <= vns_videosoc_csrbank5_core_initiator_base1_r;
	end
	if (vns_videosoc_csrbank5_core_initiator_base0_re) begin
		soc_hdmi_out0_core_initiator_csrstorage8_storage_full <= {vns_videosoc_csrbank5_core_initiator_base_backstore, vns_videosoc_csrbank5_core_initiator_base0_r};
	end
	soc_hdmi_out0_core_initiator_csrstorage8_re <= vns_videosoc_csrbank5_core_initiator_base0_re;
	if (vns_videosoc_csrbank5_core_initiator_length3_re) begin
		vns_videosoc_csrbank5_core_initiator_length_backstore[23:16] <= vns_videosoc_csrbank5_core_initiator_length3_r;
	end
	if (vns_videosoc_csrbank5_core_initiator_length2_re) begin
		vns_videosoc_csrbank5_core_initiator_length_backstore[15:8] <= vns_videosoc_csrbank5_core_initiator_length2_r;
	end
	if (vns_videosoc_csrbank5_core_initiator_length1_re) begin
		vns_videosoc_csrbank5_core_initiator_length_backstore[7:0] <= vns_videosoc_csrbank5_core_initiator_length1_r;
	end
	if (vns_videosoc_csrbank5_core_initiator_length0_re) begin
		soc_hdmi_out0_core_initiator_csrstorage9_storage_full <= {vns_videosoc_csrbank5_core_initiator_length_backstore, vns_videosoc_csrbank5_core_initiator_length0_r};
	end
	soc_hdmi_out0_core_initiator_csrstorage9_re <= vns_videosoc_csrbank5_core_initiator_length0_re;
	if (vns_videosoc_csrbank5_driver_clocking_mmcm_reset0_re) begin
		soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage_full <= vns_videosoc_csrbank5_driver_clocking_mmcm_reset0_r;
	end
	soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_re <= vns_videosoc_csrbank5_driver_clocking_mmcm_reset0_re;
	if (vns_videosoc_csrbank5_driver_clocking_mmcm_adr0_re) begin
		soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage_full[6:0] <= vns_videosoc_csrbank5_driver_clocking_mmcm_adr0_r;
	end
	soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_re <= vns_videosoc_csrbank5_driver_clocking_mmcm_adr0_re;
	if (vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w1_re) begin
		soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage_full[15:8] <= vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w1_r;
	end
	if (vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w0_re) begin
		soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage_full[7:0] <= vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w0_r;
	end
	soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_re <= vns_videosoc_csrbank5_driver_clocking_mmcm_dat_w0_re;
	vns_videosoc_interface6_bank_bus_dat_r <= 1'd0;
	if (vns_videosoc_csrbank6_sel) begin
		case (vns_videosoc_interface6_bank_bus_adr[5:0])
			1'd0: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_dna_id7_w;
			end
			1'd1: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_dna_id6_w;
			end
			2'd2: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_dna_id5_w;
			end
			2'd3: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_dna_id4_w;
			end
			3'd4: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_dna_id3_w;
			end
			3'd5: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_dna_id2_w;
			end
			3'd6: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_dna_id1_w;
			end
			3'd7: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_dna_id0_w;
			end
			4'd8: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit19_w;
			end
			4'd9: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit18_w;
			end
			4'd10: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit17_w;
			end
			4'd11: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit16_w;
			end
			4'd12: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit15_w;
			end
			4'd13: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit14_w;
			end
			4'd14: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit13_w;
			end
			4'd15: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit12_w;
			end
			5'd16: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit11_w;
			end
			5'd17: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit10_w;
			end
			5'd18: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit9_w;
			end
			5'd19: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit8_w;
			end
			5'd20: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit7_w;
			end
			5'd21: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit6_w;
			end
			5'd22: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit5_w;
			end
			5'd23: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit4_w;
			end
			5'd24: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit3_w;
			end
			5'd25: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit2_w;
			end
			5'd26: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit1_w;
			end
			5'd27: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_git_commit0_w;
			end
			5'd28: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_platform7_w;
			end
			5'd29: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_platform6_w;
			end
			5'd30: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_platform5_w;
			end
			5'd31: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_platform4_w;
			end
			6'd32: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_platform3_w;
			end
			6'd33: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_platform2_w;
			end
			6'd34: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_platform1_w;
			end
			6'd35: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_platform0_w;
			end
			6'd36: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_target7_w;
			end
			6'd37: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_target6_w;
			end
			6'd38: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_target5_w;
			end
			6'd39: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_target4_w;
			end
			6'd40: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_target3_w;
			end
			6'd41: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_target2_w;
			end
			6'd42: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_target1_w;
			end
			6'd43: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_platform_target0_w;
			end
			6'd44: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_xadc_temperature1_w;
			end
			6'd45: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_xadc_temperature0_w;
			end
			6'd46: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_xadc_vccint1_w;
			end
			6'd47: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_xadc_vccint0_w;
			end
			6'd48: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_xadc_vccaux1_w;
			end
			6'd49: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_xadc_vccaux0_w;
			end
			6'd50: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_xadc_vccbram1_w;
			end
			6'd51: begin
				vns_videosoc_interface6_bank_bus_dat_r <= vns_videosoc_csrbank6_xadc_vccbram0_w;
			end
		endcase
	end
	vns_videosoc_interface7_bank_bus_dat_r <= 1'd0;
	if (vns_videosoc_csrbank7_sel) begin
		case (vns_videosoc_interface7_bank_bus_adr[2:0])
			1'd0: begin
				vns_videosoc_interface7_bank_bus_dat_r <= soc_videosoc_oled_spimaster_ctrl_w;
			end
			1'd1: begin
				vns_videosoc_interface7_bank_bus_dat_r <= vns_videosoc_csrbank7_spi_length0_w;
			end
			2'd2: begin
				vns_videosoc_interface7_bank_bus_dat_r <= vns_videosoc_csrbank7_spi_status_w;
			end
			2'd3: begin
				vns_videosoc_interface7_bank_bus_dat_r <= vns_videosoc_csrbank7_spi_mosi0_w;
			end
			3'd4: begin
				vns_videosoc_interface7_bank_bus_dat_r <= vns_videosoc_csrbank7_gpio_out0_w;
			end
		endcase
	end
	if (vns_videosoc_csrbank7_spi_length0_re) begin
		soc_videosoc_oled_spimaster_length_storage_full[7:0] <= vns_videosoc_csrbank7_spi_length0_r;
	end
	soc_videosoc_oled_spimaster_length_re <= vns_videosoc_csrbank7_spi_length0_re;
	if (vns_videosoc_csrbank7_spi_mosi0_re) begin
		soc_videosoc_oled_spimaster_mosi_storage_full[7:0] <= vns_videosoc_csrbank7_spi_mosi0_r;
	end
	soc_videosoc_oled_spimaster_mosi_re <= vns_videosoc_csrbank7_spi_mosi0_re;
	if (vns_videosoc_csrbank7_gpio_out0_re) begin
		soc_videosoc_oled_storage_full[3:0] <= vns_videosoc_csrbank7_gpio_out0_r;
	end
	soc_videosoc_oled_re <= vns_videosoc_csrbank7_gpio_out0_re;
	vns_videosoc_interface8_bank_bus_dat_r <= 1'd0;
	if (vns_videosoc_csrbank8_sel) begin
		case (vns_videosoc_interface8_bank_bus_adr[5:0])
			1'd0: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_control0_w;
			end
			1'd1: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi0_command0_w;
			end
			2'd2: begin
				vns_videosoc_interface8_bank_bus_dat_r <= soc_videosoc_sdram_phaseinjector0_command_issue_w;
			end
			2'd3: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi0_address1_w;
			end
			3'd4: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi0_address0_w;
			end
			3'd5: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi0_baddress0_w;
			end
			3'd6: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi0_wrdata3_w;
			end
			3'd7: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi0_wrdata2_w;
			end
			4'd8: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi0_wrdata1_w;
			end
			4'd9: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi0_wrdata0_w;
			end
			4'd10: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi0_rddata3_w;
			end
			4'd11: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi0_rddata2_w;
			end
			4'd12: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi0_rddata1_w;
			end
			4'd13: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi0_rddata0_w;
			end
			4'd14: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi1_command0_w;
			end
			4'd15: begin
				vns_videosoc_interface8_bank_bus_dat_r <= soc_videosoc_sdram_phaseinjector1_command_issue_w;
			end
			5'd16: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi1_address1_w;
			end
			5'd17: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi1_address0_w;
			end
			5'd18: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi1_baddress0_w;
			end
			5'd19: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi1_wrdata3_w;
			end
			5'd20: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi1_wrdata2_w;
			end
			5'd21: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi1_wrdata1_w;
			end
			5'd22: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi1_wrdata0_w;
			end
			5'd23: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi1_rddata3_w;
			end
			5'd24: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi1_rddata2_w;
			end
			5'd25: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi1_rddata1_w;
			end
			5'd26: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi1_rddata0_w;
			end
			5'd27: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi2_command0_w;
			end
			5'd28: begin
				vns_videosoc_interface8_bank_bus_dat_r <= soc_videosoc_sdram_phaseinjector2_command_issue_w;
			end
			5'd29: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi2_address1_w;
			end
			5'd30: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi2_address0_w;
			end
			5'd31: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi2_baddress0_w;
			end
			6'd32: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi2_wrdata3_w;
			end
			6'd33: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi2_wrdata2_w;
			end
			6'd34: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi2_wrdata1_w;
			end
			6'd35: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi2_wrdata0_w;
			end
			6'd36: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi2_rddata3_w;
			end
			6'd37: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi2_rddata2_w;
			end
			6'd38: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi2_rddata1_w;
			end
			6'd39: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi2_rddata0_w;
			end
			6'd40: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi3_command0_w;
			end
			6'd41: begin
				vns_videosoc_interface8_bank_bus_dat_r <= soc_videosoc_sdram_phaseinjector3_command_issue_w;
			end
			6'd42: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi3_address1_w;
			end
			6'd43: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi3_address0_w;
			end
			6'd44: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi3_baddress0_w;
			end
			6'd45: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi3_wrdata3_w;
			end
			6'd46: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi3_wrdata2_w;
			end
			6'd47: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi3_wrdata1_w;
			end
			6'd48: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi3_wrdata0_w;
			end
			6'd49: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi3_rddata3_w;
			end
			6'd50: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi3_rddata2_w;
			end
			6'd51: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi3_rddata1_w;
			end
			6'd52: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_dfii_pi3_rddata0_w;
			end
			6'd53: begin
				vns_videosoc_interface8_bank_bus_dat_r <= soc_videosoc_sdram_bandwidth_update_w;
			end
			6'd54: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_controller_bandwidth_nreads2_w;
			end
			6'd55: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_controller_bandwidth_nreads1_w;
			end
			6'd56: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_controller_bandwidth_nreads0_w;
			end
			6'd57: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_controller_bandwidth_nwrites2_w;
			end
			6'd58: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_controller_bandwidth_nwrites1_w;
			end
			6'd59: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_controller_bandwidth_nwrites0_w;
			end
			6'd60: begin
				vns_videosoc_interface8_bank_bus_dat_r <= vns_videosoc_csrbank8_controller_bandwidth_data_width_w;
			end
		endcase
	end
	if (vns_videosoc_csrbank8_dfii_control0_re) begin
		soc_videosoc_sdram_storage_full[3:0] <= vns_videosoc_csrbank8_dfii_control0_r;
	end
	soc_videosoc_sdram_re <= vns_videosoc_csrbank8_dfii_control0_re;
	if (vns_videosoc_csrbank8_dfii_pi0_command0_re) begin
		soc_videosoc_sdram_phaseinjector0_command_storage_full[5:0] <= vns_videosoc_csrbank8_dfii_pi0_command0_r;
	end
	soc_videosoc_sdram_phaseinjector0_command_re <= vns_videosoc_csrbank8_dfii_pi0_command0_re;
	if (vns_videosoc_csrbank8_dfii_pi0_address1_re) begin
		soc_videosoc_sdram_phaseinjector0_address_storage_full[14:8] <= vns_videosoc_csrbank8_dfii_pi0_address1_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi0_address0_re) begin
		soc_videosoc_sdram_phaseinjector0_address_storage_full[7:0] <= vns_videosoc_csrbank8_dfii_pi0_address0_r;
	end
	soc_videosoc_sdram_phaseinjector0_address_re <= vns_videosoc_csrbank8_dfii_pi0_address0_re;
	if (vns_videosoc_csrbank8_dfii_pi0_baddress0_re) begin
		soc_videosoc_sdram_phaseinjector0_baddress_storage_full[2:0] <= vns_videosoc_csrbank8_dfii_pi0_baddress0_r;
	end
	soc_videosoc_sdram_phaseinjector0_baddress_re <= vns_videosoc_csrbank8_dfii_pi0_baddress0_re;
	if (vns_videosoc_csrbank8_dfii_pi0_wrdata3_re) begin
		soc_videosoc_sdram_phaseinjector0_wrdata_storage_full[31:24] <= vns_videosoc_csrbank8_dfii_pi0_wrdata3_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi0_wrdata2_re) begin
		soc_videosoc_sdram_phaseinjector0_wrdata_storage_full[23:16] <= vns_videosoc_csrbank8_dfii_pi0_wrdata2_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi0_wrdata1_re) begin
		soc_videosoc_sdram_phaseinjector0_wrdata_storage_full[15:8] <= vns_videosoc_csrbank8_dfii_pi0_wrdata1_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi0_wrdata0_re) begin
		soc_videosoc_sdram_phaseinjector0_wrdata_storage_full[7:0] <= vns_videosoc_csrbank8_dfii_pi0_wrdata0_r;
	end
	soc_videosoc_sdram_phaseinjector0_wrdata_re <= vns_videosoc_csrbank8_dfii_pi0_wrdata0_re;
	if (vns_videosoc_csrbank8_dfii_pi1_command0_re) begin
		soc_videosoc_sdram_phaseinjector1_command_storage_full[5:0] <= vns_videosoc_csrbank8_dfii_pi1_command0_r;
	end
	soc_videosoc_sdram_phaseinjector1_command_re <= vns_videosoc_csrbank8_dfii_pi1_command0_re;
	if (vns_videosoc_csrbank8_dfii_pi1_address1_re) begin
		soc_videosoc_sdram_phaseinjector1_address_storage_full[14:8] <= vns_videosoc_csrbank8_dfii_pi1_address1_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi1_address0_re) begin
		soc_videosoc_sdram_phaseinjector1_address_storage_full[7:0] <= vns_videosoc_csrbank8_dfii_pi1_address0_r;
	end
	soc_videosoc_sdram_phaseinjector1_address_re <= vns_videosoc_csrbank8_dfii_pi1_address0_re;
	if (vns_videosoc_csrbank8_dfii_pi1_baddress0_re) begin
		soc_videosoc_sdram_phaseinjector1_baddress_storage_full[2:0] <= vns_videosoc_csrbank8_dfii_pi1_baddress0_r;
	end
	soc_videosoc_sdram_phaseinjector1_baddress_re <= vns_videosoc_csrbank8_dfii_pi1_baddress0_re;
	if (vns_videosoc_csrbank8_dfii_pi1_wrdata3_re) begin
		soc_videosoc_sdram_phaseinjector1_wrdata_storage_full[31:24] <= vns_videosoc_csrbank8_dfii_pi1_wrdata3_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi1_wrdata2_re) begin
		soc_videosoc_sdram_phaseinjector1_wrdata_storage_full[23:16] <= vns_videosoc_csrbank8_dfii_pi1_wrdata2_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi1_wrdata1_re) begin
		soc_videosoc_sdram_phaseinjector1_wrdata_storage_full[15:8] <= vns_videosoc_csrbank8_dfii_pi1_wrdata1_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi1_wrdata0_re) begin
		soc_videosoc_sdram_phaseinjector1_wrdata_storage_full[7:0] <= vns_videosoc_csrbank8_dfii_pi1_wrdata0_r;
	end
	soc_videosoc_sdram_phaseinjector1_wrdata_re <= vns_videosoc_csrbank8_dfii_pi1_wrdata0_re;
	if (vns_videosoc_csrbank8_dfii_pi2_command0_re) begin
		soc_videosoc_sdram_phaseinjector2_command_storage_full[5:0] <= vns_videosoc_csrbank8_dfii_pi2_command0_r;
	end
	soc_videosoc_sdram_phaseinjector2_command_re <= vns_videosoc_csrbank8_dfii_pi2_command0_re;
	if (vns_videosoc_csrbank8_dfii_pi2_address1_re) begin
		soc_videosoc_sdram_phaseinjector2_address_storage_full[14:8] <= vns_videosoc_csrbank8_dfii_pi2_address1_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi2_address0_re) begin
		soc_videosoc_sdram_phaseinjector2_address_storage_full[7:0] <= vns_videosoc_csrbank8_dfii_pi2_address0_r;
	end
	soc_videosoc_sdram_phaseinjector2_address_re <= vns_videosoc_csrbank8_dfii_pi2_address0_re;
	if (vns_videosoc_csrbank8_dfii_pi2_baddress0_re) begin
		soc_videosoc_sdram_phaseinjector2_baddress_storage_full[2:0] <= vns_videosoc_csrbank8_dfii_pi2_baddress0_r;
	end
	soc_videosoc_sdram_phaseinjector2_baddress_re <= vns_videosoc_csrbank8_dfii_pi2_baddress0_re;
	if (vns_videosoc_csrbank8_dfii_pi2_wrdata3_re) begin
		soc_videosoc_sdram_phaseinjector2_wrdata_storage_full[31:24] <= vns_videosoc_csrbank8_dfii_pi2_wrdata3_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi2_wrdata2_re) begin
		soc_videosoc_sdram_phaseinjector2_wrdata_storage_full[23:16] <= vns_videosoc_csrbank8_dfii_pi2_wrdata2_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi2_wrdata1_re) begin
		soc_videosoc_sdram_phaseinjector2_wrdata_storage_full[15:8] <= vns_videosoc_csrbank8_dfii_pi2_wrdata1_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi2_wrdata0_re) begin
		soc_videosoc_sdram_phaseinjector2_wrdata_storage_full[7:0] <= vns_videosoc_csrbank8_dfii_pi2_wrdata0_r;
	end
	soc_videosoc_sdram_phaseinjector2_wrdata_re <= vns_videosoc_csrbank8_dfii_pi2_wrdata0_re;
	if (vns_videosoc_csrbank8_dfii_pi3_command0_re) begin
		soc_videosoc_sdram_phaseinjector3_command_storage_full[5:0] <= vns_videosoc_csrbank8_dfii_pi3_command0_r;
	end
	soc_videosoc_sdram_phaseinjector3_command_re <= vns_videosoc_csrbank8_dfii_pi3_command0_re;
	if (vns_videosoc_csrbank8_dfii_pi3_address1_re) begin
		soc_videosoc_sdram_phaseinjector3_address_storage_full[14:8] <= vns_videosoc_csrbank8_dfii_pi3_address1_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi3_address0_re) begin
		soc_videosoc_sdram_phaseinjector3_address_storage_full[7:0] <= vns_videosoc_csrbank8_dfii_pi3_address0_r;
	end
	soc_videosoc_sdram_phaseinjector3_address_re <= vns_videosoc_csrbank8_dfii_pi3_address0_re;
	if (vns_videosoc_csrbank8_dfii_pi3_baddress0_re) begin
		soc_videosoc_sdram_phaseinjector3_baddress_storage_full[2:0] <= vns_videosoc_csrbank8_dfii_pi3_baddress0_r;
	end
	soc_videosoc_sdram_phaseinjector3_baddress_re <= vns_videosoc_csrbank8_dfii_pi3_baddress0_re;
	if (vns_videosoc_csrbank8_dfii_pi3_wrdata3_re) begin
		soc_videosoc_sdram_phaseinjector3_wrdata_storage_full[31:24] <= vns_videosoc_csrbank8_dfii_pi3_wrdata3_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi3_wrdata2_re) begin
		soc_videosoc_sdram_phaseinjector3_wrdata_storage_full[23:16] <= vns_videosoc_csrbank8_dfii_pi3_wrdata2_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi3_wrdata1_re) begin
		soc_videosoc_sdram_phaseinjector3_wrdata_storage_full[15:8] <= vns_videosoc_csrbank8_dfii_pi3_wrdata1_r;
	end
	if (vns_videosoc_csrbank8_dfii_pi3_wrdata0_re) begin
		soc_videosoc_sdram_phaseinjector3_wrdata_storage_full[7:0] <= vns_videosoc_csrbank8_dfii_pi3_wrdata0_r;
	end
	soc_videosoc_sdram_phaseinjector3_wrdata_re <= vns_videosoc_csrbank8_dfii_pi3_wrdata0_re;
	vns_videosoc_interface9_bank_bus_dat_r <= 1'd0;
	if (vns_videosoc_csrbank9_sel) begin
		case (vns_videosoc_interface9_bank_bus_adr[1:0])
			1'd0: begin
				vns_videosoc_interface9_bank_bus_dat_r <= vns_videosoc_csrbank9_bitbang0_w;
			end
			1'd1: begin
				vns_videosoc_interface9_bank_bus_dat_r <= vns_videosoc_csrbank9_miso_w;
			end
			2'd2: begin
				vns_videosoc_interface9_bank_bus_dat_r <= vns_videosoc_csrbank9_bitbang_en0_w;
			end
		endcase
	end
	if (vns_videosoc_csrbank9_bitbang0_re) begin
		soc_videosoc_bitbang_storage_full[3:0] <= vns_videosoc_csrbank9_bitbang0_r;
	end
	soc_videosoc_bitbang_re <= vns_videosoc_csrbank9_bitbang0_re;
	if (vns_videosoc_csrbank9_bitbang_en0_re) begin
		soc_videosoc_bitbang_en_storage_full <= vns_videosoc_csrbank9_bitbang_en0_r;
	end
	soc_videosoc_bitbang_en_re <= vns_videosoc_csrbank9_bitbang_en0_re;
	vns_videosoc_interface10_bank_bus_dat_r <= 1'd0;
	if (vns_videosoc_csrbank10_sel) begin
		case (vns_videosoc_interface10_bank_bus_adr[4:0])
			1'd0: begin
				vns_videosoc_interface10_bank_bus_dat_r <= vns_videosoc_csrbank10_load3_w;
			end
			1'd1: begin
				vns_videosoc_interface10_bank_bus_dat_r <= vns_videosoc_csrbank10_load2_w;
			end
			2'd2: begin
				vns_videosoc_interface10_bank_bus_dat_r <= vns_videosoc_csrbank10_load1_w;
			end
			2'd3: begin
				vns_videosoc_interface10_bank_bus_dat_r <= vns_videosoc_csrbank10_load0_w;
			end
			3'd4: begin
				vns_videosoc_interface10_bank_bus_dat_r <= vns_videosoc_csrbank10_reload3_w;
			end
			3'd5: begin
				vns_videosoc_interface10_bank_bus_dat_r <= vns_videosoc_csrbank10_reload2_w;
			end
			3'd6: begin
				vns_videosoc_interface10_bank_bus_dat_r <= vns_videosoc_csrbank10_reload1_w;
			end
			3'd7: begin
				vns_videosoc_interface10_bank_bus_dat_r <= vns_videosoc_csrbank10_reload0_w;
			end
			4'd8: begin
				vns_videosoc_interface10_bank_bus_dat_r <= vns_videosoc_csrbank10_en0_w;
			end
			4'd9: begin
				vns_videosoc_interface10_bank_bus_dat_r <= soc_videosoc_videosoc_update_value_w;
			end
			4'd10: begin
				vns_videosoc_interface10_bank_bus_dat_r <= vns_videosoc_csrbank10_value3_w;
			end
			4'd11: begin
				vns_videosoc_interface10_bank_bus_dat_r <= vns_videosoc_csrbank10_value2_w;
			end
			4'd12: begin
				vns_videosoc_interface10_bank_bus_dat_r <= vns_videosoc_csrbank10_value1_w;
			end
			4'd13: begin
				vns_videosoc_interface10_bank_bus_dat_r <= vns_videosoc_csrbank10_value0_w;
			end
			4'd14: begin
				vns_videosoc_interface10_bank_bus_dat_r <= soc_videosoc_videosoc_eventmanager_status_w;
			end
			4'd15: begin
				vns_videosoc_interface10_bank_bus_dat_r <= soc_videosoc_videosoc_eventmanager_pending_w;
			end
			5'd16: begin
				vns_videosoc_interface10_bank_bus_dat_r <= vns_videosoc_csrbank10_ev_enable0_w;
			end
		endcase
	end
	if (vns_videosoc_csrbank10_load3_re) begin
		soc_videosoc_videosoc_load_storage_full[31:24] <= vns_videosoc_csrbank10_load3_r;
	end
	if (vns_videosoc_csrbank10_load2_re) begin
		soc_videosoc_videosoc_load_storage_full[23:16] <= vns_videosoc_csrbank10_load2_r;
	end
	if (vns_videosoc_csrbank10_load1_re) begin
		soc_videosoc_videosoc_load_storage_full[15:8] <= vns_videosoc_csrbank10_load1_r;
	end
	if (vns_videosoc_csrbank10_load0_re) begin
		soc_videosoc_videosoc_load_storage_full[7:0] <= vns_videosoc_csrbank10_load0_r;
	end
	soc_videosoc_videosoc_load_re <= vns_videosoc_csrbank10_load0_re;
	if (vns_videosoc_csrbank10_reload3_re) begin
		soc_videosoc_videosoc_reload_storage_full[31:24] <= vns_videosoc_csrbank10_reload3_r;
	end
	if (vns_videosoc_csrbank10_reload2_re) begin
		soc_videosoc_videosoc_reload_storage_full[23:16] <= vns_videosoc_csrbank10_reload2_r;
	end
	if (vns_videosoc_csrbank10_reload1_re) begin
		soc_videosoc_videosoc_reload_storage_full[15:8] <= vns_videosoc_csrbank10_reload1_r;
	end
	if (vns_videosoc_csrbank10_reload0_re) begin
		soc_videosoc_videosoc_reload_storage_full[7:0] <= vns_videosoc_csrbank10_reload0_r;
	end
	soc_videosoc_videosoc_reload_re <= vns_videosoc_csrbank10_reload0_re;
	if (vns_videosoc_csrbank10_en0_re) begin
		soc_videosoc_videosoc_en_storage_full <= vns_videosoc_csrbank10_en0_r;
	end
	soc_videosoc_videosoc_en_re <= vns_videosoc_csrbank10_en0_re;
	if (vns_videosoc_csrbank10_ev_enable0_re) begin
		soc_videosoc_videosoc_eventmanager_storage_full <= vns_videosoc_csrbank10_ev_enable0_r;
	end
	soc_videosoc_videosoc_eventmanager_re <= vns_videosoc_csrbank10_ev_enable0_re;
	vns_videosoc_interface11_bank_bus_dat_r <= 1'd0;
	if (vns_videosoc_csrbank11_sel) begin
		case (vns_videosoc_interface11_bank_bus_adr[2:0])
			1'd0: begin
				vns_videosoc_interface11_bank_bus_dat_r <= soc_videosoc_uart_rxtx_w;
			end
			1'd1: begin
				vns_videosoc_interface11_bank_bus_dat_r <= vns_videosoc_csrbank11_txfull_w;
			end
			2'd2: begin
				vns_videosoc_interface11_bank_bus_dat_r <= vns_videosoc_csrbank11_rxempty_w;
			end
			2'd3: begin
				vns_videosoc_interface11_bank_bus_dat_r <= soc_videosoc_uart_status_w;
			end
			3'd4: begin
				vns_videosoc_interface11_bank_bus_dat_r <= soc_videosoc_uart_pending_w;
			end
			3'd5: begin
				vns_videosoc_interface11_bank_bus_dat_r <= vns_videosoc_csrbank11_ev_enable0_w;
			end
		endcase
	end
	if (vns_videosoc_csrbank11_ev_enable0_re) begin
		soc_videosoc_uart_storage_full[1:0] <= vns_videosoc_csrbank11_ev_enable0_r;
	end
	soc_videosoc_uart_re <= vns_videosoc_csrbank11_ev_enable0_re;
	vns_videosoc_interface12_bank_bus_dat_r <= 1'd0;
	if (vns_videosoc_csrbank12_sel) begin
		case (vns_videosoc_interface12_bank_bus_adr[1:0])
			1'd0: begin
				vns_videosoc_interface12_bank_bus_dat_r <= vns_videosoc_csrbank12_tuning_word3_w;
			end
			1'd1: begin
				vns_videosoc_interface12_bank_bus_dat_r <= vns_videosoc_csrbank12_tuning_word2_w;
			end
			2'd2: begin
				vns_videosoc_interface12_bank_bus_dat_r <= vns_videosoc_csrbank12_tuning_word1_w;
			end
			2'd3: begin
				vns_videosoc_interface12_bank_bus_dat_r <= vns_videosoc_csrbank12_tuning_word0_w;
			end
		endcase
	end
	if (vns_videosoc_csrbank12_tuning_word3_re) begin
		soc_videosoc_uart_phy_storage_full[31:24] <= vns_videosoc_csrbank12_tuning_word3_r;
	end
	if (vns_videosoc_csrbank12_tuning_word2_re) begin
		soc_videosoc_uart_phy_storage_full[23:16] <= vns_videosoc_csrbank12_tuning_word2_r;
	end
	if (vns_videosoc_csrbank12_tuning_word1_re) begin
		soc_videosoc_uart_phy_storage_full[15:8] <= vns_videosoc_csrbank12_tuning_word1_r;
	end
	if (vns_videosoc_csrbank12_tuning_word0_re) begin
		soc_videosoc_uart_phy_storage_full[7:0] <= vns_videosoc_csrbank12_tuning_word0_r;
	end
	soc_videosoc_uart_phy_re <= vns_videosoc_csrbank12_tuning_word0_re;
	if (sys_rst) begin
		soc_videosoc_videosoc_rom_bus_ack <= 1'd0;
		soc_videosoc_videosoc_sram_bus_ack <= 1'd0;
		soc_videosoc_videosoc_interface_adr <= 14'd0;
		soc_videosoc_videosoc_interface_we <= 1'd0;
		soc_videosoc_videosoc_interface_dat_w <= 8'd0;
		soc_videosoc_videosoc_bus_wishbone_dat_r <= 32'd0;
		soc_videosoc_videosoc_bus_wishbone_ack <= 1'd0;
		soc_videosoc_videosoc_counter <= 2'd0;
		soc_videosoc_videosoc_load_storage_full <= 32'd0;
		soc_videosoc_videosoc_load_re <= 1'd0;
		soc_videosoc_videosoc_reload_storage_full <= 32'd0;
		soc_videosoc_videosoc_reload_re <= 1'd0;
		soc_videosoc_videosoc_en_storage_full <= 1'd0;
		soc_videosoc_videosoc_en_re <= 1'd0;
		soc_videosoc_videosoc_value_status <= 32'd0;
		soc_videosoc_videosoc_zero_pending <= 1'd0;
		soc_videosoc_videosoc_zero_old_trigger <= 1'd0;
		soc_videosoc_videosoc_eventmanager_storage_full <= 1'd0;
		soc_videosoc_videosoc_eventmanager_re <= 1'd0;
		soc_videosoc_videosoc_value <= 32'd0;
		soc_videosoc_uart_tx_pending <= 1'd0;
		soc_videosoc_uart_tx_old_trigger <= 1'd0;
		soc_videosoc_uart_rx_pending <= 1'd0;
		soc_videosoc_uart_rx_old_trigger <= 1'd0;
		soc_videosoc_uart_storage_full <= 2'd0;
		soc_videosoc_uart_re <= 1'd0;
		soc_videosoc_uart_tx_fifo_level <= 5'd0;
		soc_videosoc_uart_tx_fifo_produce <= 4'd0;
		soc_videosoc_uart_tx_fifo_consume <= 4'd0;
		soc_videosoc_uart_rx_fifo_level <= 5'd0;
		soc_videosoc_uart_rx_fifo_produce <= 4'd0;
		soc_videosoc_uart_rx_fifo_consume <= 4'd0;
		soc_videosoc_bridge_count <= 24'd10000000;
		serial_tx <= 1'd1;
		soc_videosoc_uart_phy_storage_full <= 32'd4947802;
		soc_videosoc_uart_phy_re <= 1'd0;
		soc_videosoc_uart_phy_sink_ready <= 1'd0;
		soc_videosoc_uart_phy_uart_clk_txen <= 1'd0;
		soc_videosoc_uart_phy_phase_accumulator_tx <= 32'd0;
		soc_videosoc_uart_phy_tx_reg <= 8'd0;
		soc_videosoc_uart_phy_tx_bitcount <= 4'd0;
		soc_videosoc_uart_phy_tx_busy <= 1'd0;
		soc_videosoc_uart_phy_source_valid <= 1'd0;
		soc_videosoc_uart_phy_uart_clk_rxen <= 1'd0;
		soc_videosoc_uart_phy_phase_accumulator_rx <= 32'd0;
		soc_videosoc_uart_phy_rx_r <= 1'd0;
		soc_videosoc_uart_phy_rx_reg <= 8'd0;
		soc_videosoc_uart_phy_rx_bitcount <= 4'd0;
		soc_videosoc_uart_phy_rx_busy <= 1'd0;
		soc_videosoc_info_dna_status <= 57'd0;
		soc_videosoc_info_dna_cnt <= 7'd0;
		soc_videosoc_info_temperature_status <= 12'd0;
		soc_videosoc_info_vccint_status <= 12'd0;
		soc_videosoc_info_vccaux_status <= 12'd0;
		soc_videosoc_info_vccbram_status <= 12'd0;
		soc_videosoc_oled_spi_pads_clk <= 1'd0;
		soc_videosoc_oled_spi_pads_mosi <= 1'd0;
		soc_videosoc_oled_spimaster_length_storage_full <= 8'd0;
		soc_videosoc_oled_spimaster_length_re <= 1'd0;
		soc_videosoc_oled_spimaster_mosi_storage_full <= 8'd0;
		soc_videosoc_oled_spimaster_mosi_re <= 1'd0;
		soc_videosoc_oled_spimaster_i <= 4'd0;
		soc_videosoc_oled_spimaster_cnt <= 8'd0;
		soc_videosoc_oled_spimaster_sr_mosi <= 8'd0;
		soc_videosoc_oled_storage_full <= 4'd0;
		soc_videosoc_oled_re <= 1'd0;
		soc_videosoc_ddrphy_storage_full <= 2'd0;
		soc_videosoc_ddrphy_re <= 1'd0;
		soc_videosoc_ddrphy_dfi_p0_rddata_valid <= 1'd0;
		soc_videosoc_ddrphy_dfi_p1_rddata_valid <= 1'd0;
		soc_videosoc_ddrphy_dfi_p2_rddata_valid <= 1'd0;
		soc_videosoc_ddrphy_dfi_p3_rddata_valid <= 1'd0;
		soc_videosoc_ddrphy_oe_dqs <= 1'd0;
		soc_videosoc_ddrphy_oe_dq <= 1'd0;
		soc_videosoc_ddrphy_n_rddata_en0 <= 1'd0;
		soc_videosoc_ddrphy_n_rddata_en1 <= 1'd0;
		soc_videosoc_ddrphy_n_rddata_en2 <= 1'd0;
		soc_videosoc_ddrphy_n_rddata_en3 <= 1'd0;
		soc_videosoc_ddrphy_n_rddata_en4 <= 1'd0;
		soc_videosoc_ddrphy_last_wrdata_en <= 4'd0;
		soc_videosoc_sdram_storage_full <= 4'd0;
		soc_videosoc_sdram_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector0_command_storage_full <= 6'd0;
		soc_videosoc_sdram_phaseinjector0_command_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector0_address_storage_full <= 15'd0;
		soc_videosoc_sdram_phaseinjector0_address_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector0_baddress_storage_full <= 3'd0;
		soc_videosoc_sdram_phaseinjector0_baddress_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector0_wrdata_storage_full <= 32'd0;
		soc_videosoc_sdram_phaseinjector0_wrdata_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector0_status <= 32'd0;
		soc_videosoc_sdram_phaseinjector1_command_storage_full <= 6'd0;
		soc_videosoc_sdram_phaseinjector1_command_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector1_address_storage_full <= 15'd0;
		soc_videosoc_sdram_phaseinjector1_address_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector1_baddress_storage_full <= 3'd0;
		soc_videosoc_sdram_phaseinjector1_baddress_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector1_wrdata_storage_full <= 32'd0;
		soc_videosoc_sdram_phaseinjector1_wrdata_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector1_status <= 32'd0;
		soc_videosoc_sdram_phaseinjector2_command_storage_full <= 6'd0;
		soc_videosoc_sdram_phaseinjector2_command_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector2_address_storage_full <= 15'd0;
		soc_videosoc_sdram_phaseinjector2_address_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector2_baddress_storage_full <= 3'd0;
		soc_videosoc_sdram_phaseinjector2_baddress_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector2_wrdata_storage_full <= 32'd0;
		soc_videosoc_sdram_phaseinjector2_wrdata_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector2_status <= 32'd0;
		soc_videosoc_sdram_phaseinjector3_command_storage_full <= 6'd0;
		soc_videosoc_sdram_phaseinjector3_command_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector3_address_storage_full <= 15'd0;
		soc_videosoc_sdram_phaseinjector3_address_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector3_baddress_storage_full <= 3'd0;
		soc_videosoc_sdram_phaseinjector3_baddress_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector3_wrdata_storage_full <= 32'd0;
		soc_videosoc_sdram_phaseinjector3_wrdata_re <= 1'd0;
		soc_videosoc_sdram_phaseinjector3_status <= 32'd0;
		soc_videosoc_sdram_dfi_p0_cas_n <= 1'd1;
		soc_videosoc_sdram_dfi_p0_ras_n <= 1'd1;
		soc_videosoc_sdram_dfi_p0_we_n <= 1'd1;
		soc_videosoc_sdram_dfi_p0_wrdata_en <= 1'd0;
		soc_videosoc_sdram_dfi_p0_rddata_en <= 1'd0;
		soc_videosoc_sdram_dfi_p1_cas_n <= 1'd1;
		soc_videosoc_sdram_dfi_p1_ras_n <= 1'd1;
		soc_videosoc_sdram_dfi_p1_we_n <= 1'd1;
		soc_videosoc_sdram_dfi_p1_wrdata_en <= 1'd0;
		soc_videosoc_sdram_dfi_p1_rddata_en <= 1'd0;
		soc_videosoc_sdram_dfi_p2_cas_n <= 1'd1;
		soc_videosoc_sdram_dfi_p2_ras_n <= 1'd1;
		soc_videosoc_sdram_dfi_p2_we_n <= 1'd1;
		soc_videosoc_sdram_dfi_p2_wrdata_en <= 1'd0;
		soc_videosoc_sdram_dfi_p2_rddata_en <= 1'd0;
		soc_videosoc_sdram_dfi_p3_cas_n <= 1'd1;
		soc_videosoc_sdram_dfi_p3_ras_n <= 1'd1;
		soc_videosoc_sdram_dfi_p3_we_n <= 1'd1;
		soc_videosoc_sdram_dfi_p3_wrdata_en <= 1'd0;
		soc_videosoc_sdram_dfi_p3_rddata_en <= 1'd0;
		soc_videosoc_sdram_seq_done <= 1'd0;
		soc_videosoc_sdram_counter <= 5'd0;
		soc_videosoc_sdram_count <= 10'd782;
		soc_videosoc_sdram_bankmachine0_level <= 4'd0;
		soc_videosoc_sdram_bankmachine0_produce <= 3'd0;
		soc_videosoc_sdram_bankmachine0_consume <= 3'd0;
		soc_videosoc_sdram_bankmachine0_has_openrow <= 1'd0;
		soc_videosoc_sdram_bankmachine0_count <= 3'd5;
		soc_videosoc_sdram_bankmachine1_level <= 4'd0;
		soc_videosoc_sdram_bankmachine1_produce <= 3'd0;
		soc_videosoc_sdram_bankmachine1_consume <= 3'd0;
		soc_videosoc_sdram_bankmachine1_has_openrow <= 1'd0;
		soc_videosoc_sdram_bankmachine1_count <= 3'd5;
		soc_videosoc_sdram_bankmachine2_level <= 4'd0;
		soc_videosoc_sdram_bankmachine2_produce <= 3'd0;
		soc_videosoc_sdram_bankmachine2_consume <= 3'd0;
		soc_videosoc_sdram_bankmachine2_has_openrow <= 1'd0;
		soc_videosoc_sdram_bankmachine2_count <= 3'd5;
		soc_videosoc_sdram_bankmachine3_level <= 4'd0;
		soc_videosoc_sdram_bankmachine3_produce <= 3'd0;
		soc_videosoc_sdram_bankmachine3_consume <= 3'd0;
		soc_videosoc_sdram_bankmachine3_has_openrow <= 1'd0;
		soc_videosoc_sdram_bankmachine3_count <= 3'd5;
		soc_videosoc_sdram_bankmachine4_level <= 4'd0;
		soc_videosoc_sdram_bankmachine4_produce <= 3'd0;
		soc_videosoc_sdram_bankmachine4_consume <= 3'd0;
		soc_videosoc_sdram_bankmachine4_has_openrow <= 1'd0;
		soc_videosoc_sdram_bankmachine4_count <= 3'd5;
		soc_videosoc_sdram_bankmachine5_level <= 4'd0;
		soc_videosoc_sdram_bankmachine5_produce <= 3'd0;
		soc_videosoc_sdram_bankmachine5_consume <= 3'd0;
		soc_videosoc_sdram_bankmachine5_has_openrow <= 1'd0;
		soc_videosoc_sdram_bankmachine5_count <= 3'd5;
		soc_videosoc_sdram_bankmachine6_level <= 4'd0;
		soc_videosoc_sdram_bankmachine6_produce <= 3'd0;
		soc_videosoc_sdram_bankmachine6_consume <= 3'd0;
		soc_videosoc_sdram_bankmachine6_has_openrow <= 1'd0;
		soc_videosoc_sdram_bankmachine6_count <= 3'd5;
		soc_videosoc_sdram_bankmachine7_level <= 4'd0;
		soc_videosoc_sdram_bankmachine7_produce <= 3'd0;
		soc_videosoc_sdram_bankmachine7_consume <= 3'd0;
		soc_videosoc_sdram_bankmachine7_has_openrow <= 1'd0;
		soc_videosoc_sdram_bankmachine7_count <= 3'd5;
		soc_videosoc_sdram_choose_cmd_grant <= 3'd0;
		soc_videosoc_sdram_choose_req_grant <= 3'd0;
		soc_videosoc_sdram_time0 <= 5'd0;
		soc_videosoc_sdram_time1 <= 4'd0;
		soc_videosoc_sdram_bandwidth_nreads_status <= 24'd0;
		soc_videosoc_sdram_bandwidth_nwrites_status <= 24'd0;
		soc_videosoc_sdram_bandwidth_cmd_valid <= 1'd0;
		soc_videosoc_sdram_bandwidth_cmd_ready <= 1'd0;
		soc_videosoc_sdram_bandwidth_cmd_is_read <= 1'd0;
		soc_videosoc_sdram_bandwidth_cmd_is_write <= 1'd0;
		soc_videosoc_sdram_bandwidth_counter <= 24'd0;
		soc_videosoc_sdram_bandwidth_period <= 1'd0;
		soc_videosoc_sdram_bandwidth_nreads <= 24'd0;
		soc_videosoc_sdram_bandwidth_nwrites <= 24'd0;
		soc_videosoc_sdram_bandwidth_nreads_r <= 24'd0;
		soc_videosoc_sdram_bandwidth_nwrites_r <= 24'd0;
		soc_videosoc_adr_offset_r <= 2'd0;
		soc_videosoc_bus_ack <= 1'd0;
		soc_videosoc_bitbang_storage_full <= 4'd0;
		soc_videosoc_bitbang_re <= 1'd0;
		soc_videosoc_bitbang_en_storage_full <= 1'd0;
		soc_videosoc_bitbang_en_re <= 1'd0;
		soc_videosoc_cs_n <= 1'd1;
		soc_videosoc_clk1 <= 1'd0;
		soc_videosoc_sr <= 32'd0;
		soc_videosoc_i <= 1'd0;
		soc_videosoc_miso <= 1'd0;
		soc_videosoc_counter <= 8'd0;
		soc_ethphy_reset_storage_full <= 1'd0;
		soc_ethphy_reset_re <= 1'd0;
		soc_ethphy_counter <= 9'd0;
		soc_ethphy_storage_full <= 3'd0;
		soc_ethphy_re <= 1'd0;
		soc_ethmac_tx_cdc_graycounter0_q <= 7'd0;
		soc_ethmac_tx_cdc_graycounter0_q_binary <= 7'd0;
		soc_ethmac_rx_cdc_graycounter1_q <= 7'd0;
		soc_ethmac_rx_cdc_graycounter1_q_binary <= 7'd0;
		soc_ethmac_writer_storage_full <= 1'd0;
		soc_ethmac_writer_re <= 1'd0;
		soc_ethmac_writer_counter <= 32'd0;
		soc_ethmac_writer_slot <= 1'd0;
		soc_ethmac_writer_fifo_level <= 2'd0;
		soc_ethmac_writer_fifo_produce <= 1'd0;
		soc_ethmac_writer_fifo_consume <= 1'd0;
		soc_ethmac_reader_slot_storage_full <= 1'd0;
		soc_ethmac_reader_slot_re <= 1'd0;
		soc_ethmac_reader_length_storage_full <= 11'd0;
		soc_ethmac_reader_length_re <= 1'd0;
		soc_ethmac_reader_done_pending <= 1'd0;
		soc_ethmac_reader_eventmanager_storage_full <= 1'd0;
		soc_ethmac_reader_eventmanager_re <= 1'd0;
		soc_ethmac_reader_fifo_level <= 2'd0;
		soc_ethmac_reader_fifo_produce <= 1'd0;
		soc_ethmac_reader_fifo_consume <= 1'd0;
		soc_ethmac_reader_counter <= 11'd0;
		soc_ethmac_sram0_bus_ack0 <= 1'd0;
		soc_ethmac_sram1_bus_ack0 <= 1'd0;
		soc_ethmac_sram0_bus_ack1 <= 1'd0;
		soc_ethmac_sram1_bus_ack1 <= 1'd0;
		soc_ethmac_slave_sel_r <= 4'd0;
		soc_edid_storage_full <= 1'd0;
		soc_edid_re <= 1'd0;
		soc_edid_sda_i <= 1'd0;
		soc_edid_sda_drv_reg <= 1'd0;
		soc_edid_scl_i <= 1'd0;
		soc_edid_samp_count <= 6'd0;
		soc_edid_samp_carry <= 1'd0;
		soc_edid_scl_r <= 1'd0;
		soc_edid_sda_r <= 1'd0;
		soc_edid_din <= 8'd0;
		soc_edid_counter <= 4'd0;
		soc_edid_is_read <= 1'd0;
		soc_edid_offset_counter <= 7'd0;
		soc_edid_data_bit <= 1'd0;
		soc_edid_data_drv <= 1'd0;
		soc_mmcm_reset_storage_full <= 1'd1;
		soc_mmcm_reset_re <= 1'd0;
		soc_mmcm_drdy_status <= 1'd0;
		soc_mmcm_adr_storage_full <= 7'd0;
		soc_mmcm_adr_re <= 1'd0;
		soc_mmcm_dat_w_storage_full <= 16'd0;
		soc_mmcm_dat_w_re <= 1'd0;
		soc_wer0_status <= 24'd0;
		soc_wer0_wer_counter_sys <= 24'd0;
		soc_wer1_status <= 24'd0;
		soc_wer1_wer_counter_sys <= 24'd0;
		soc_wer2_status <= 24'd0;
		soc_wer2_wer_counter_sys <= 24'd0;
		soc_frame_fifo_graycounter1_q <= 10'd0;
		soc_frame_fifo_graycounter1_q_binary <= 10'd0;
		soc_frame_overflow_mask <= 1'd0;
		soc_dma_frame_size_storage_full <= 29'd0;
		soc_dma_frame_size_re <= 1'd0;
		soc_dma_slot_array_slot0_status_storage_full <= 2'd0;
		soc_dma_slot_array_slot0_status_re <= 1'd0;
		soc_dma_slot_array_slot0_address_storage_full <= 29'd0;
		soc_dma_slot_array_slot0_address_re <= 1'd0;
		soc_dma_slot_array_slot1_status_storage_full <= 2'd0;
		soc_dma_slot_array_slot1_status_re <= 1'd0;
		soc_dma_slot_array_slot1_address_storage_full <= 29'd0;
		soc_dma_slot_array_slot1_address_re <= 1'd0;
		soc_dma_slot_array_storage_full <= 2'd0;
		soc_dma_slot_array_re <= 1'd0;
		soc_dma_slot_array_current_slot <= 1'd0;
		soc_dma_current_address <= 25'd0;
		soc_dma_mwords_remaining <= 25'd0;
		soc_dma_fifo_level <= 5'd0;
		soc_dma_fifo_produce <= 4'd0;
		soc_dma_fifo_consume <= 4'd0;
		soc_hdmi_in0_freq_period_counter <= 32'd0;
		soc_hdmi_in0_freq_sampler_o <= 32'd0;
		soc_hdmi_in0_freq_sampler_counter <= 32'd0;
		soc_hdmi_in0_freq_sampler_i_d <= 6'd0;
		soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q <= 3'd0;
		soc_hdmi_out0_dram_port_cmd_fifo_graycounter1_q_binary <= 3'd0;
		soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q <= 5'd0;
		soc_hdmi_out0_dram_port_rdata_fifo_graycounter0_q_binary <= 5'd0;
		soc_hdmi_out0_core_underflow_enable_storage_full <= 1'd0;
		soc_hdmi_out0_core_underflow_enable_re <= 1'd0;
		soc_hdmi_out0_core_initiator_cdc_graycounter0_q <= 2'd0;
		soc_hdmi_out0_core_initiator_cdc_graycounter0_q_binary <= 2'd0;
		soc_hdmi_out0_core_initiator_enable_storage_full <= 1'd0;
		soc_hdmi_out0_core_initiator_enable_re <= 1'd0;
		soc_hdmi_out0_core_initiator_csrstorage0_storage_full <= 12'd0;
		soc_hdmi_out0_core_initiator_csrstorage0_re <= 1'd0;
		soc_hdmi_out0_core_initiator_csrstorage1_storage_full <= 12'd0;
		soc_hdmi_out0_core_initiator_csrstorage1_re <= 1'd0;
		soc_hdmi_out0_core_initiator_csrstorage2_storage_full <= 12'd0;
		soc_hdmi_out0_core_initiator_csrstorage2_re <= 1'd0;
		soc_hdmi_out0_core_initiator_csrstorage3_storage_full <= 12'd0;
		soc_hdmi_out0_core_initiator_csrstorage3_re <= 1'd0;
		soc_hdmi_out0_core_initiator_csrstorage4_storage_full <= 12'd0;
		soc_hdmi_out0_core_initiator_csrstorage4_re <= 1'd0;
		soc_hdmi_out0_core_initiator_csrstorage5_storage_full <= 12'd0;
		soc_hdmi_out0_core_initiator_csrstorage5_re <= 1'd0;
		soc_hdmi_out0_core_initiator_csrstorage6_storage_full <= 12'd0;
		soc_hdmi_out0_core_initiator_csrstorage6_re <= 1'd0;
		soc_hdmi_out0_core_initiator_csrstorage7_storage_full <= 12'd0;
		soc_hdmi_out0_core_initiator_csrstorage7_re <= 1'd0;
		soc_hdmi_out0_core_initiator_csrstorage8_storage_full <= 32'd0;
		soc_hdmi_out0_core_initiator_csrstorage8_re <= 1'd0;
		soc_hdmi_out0_core_initiator_csrstorage9_storage_full <= 32'd0;
		soc_hdmi_out0_core_initiator_csrstorage9_re <= 1'd0;
		soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage_full <= 1'd0;
		soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_re <= 1'd0;
		soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy_status <= 1'd0;
		soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage_full <= 7'd0;
		soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_re <= 1'd0;
		soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage_full <= 16'd0;
		soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_re <= 1'd0;
		vns_wishbonestreamingbridge_state <= 3'd0;
		vns_oled_state <= 2'd0;
		vns_refresher_state <= 2'd0;
		vns_bankmachine0_state <= 3'd0;
		vns_bankmachine1_state <= 3'd0;
		vns_bankmachine2_state <= 3'd0;
		vns_bankmachine3_state <= 3'd0;
		vns_bankmachine4_state <= 3'd0;
		vns_bankmachine5_state <= 3'd0;
		vns_bankmachine6_state <= 3'd0;
		vns_bankmachine7_state <= 3'd0;
		vns_multiplexer_state <= 4'd0;
		vns_roundrobin0_grant <= 2'd0;
		vns_roundrobin1_grant <= 2'd0;
		vns_roundrobin2_grant <= 2'd0;
		vns_roundrobin3_grant <= 2'd0;
		vns_roundrobin4_grant <= 2'd0;
		vns_roundrobin5_grant <= 2'd0;
		vns_roundrobin6_grant <= 2'd0;
		vns_roundrobin7_grant <= 2'd0;
		vns_new_master_wdata_ready0 <= 1'd0;
		vns_new_master_wdata_ready1 <= 1'd0;
		vns_new_master_wdata_ready2 <= 1'd0;
		vns_new_master_wdata_ready3 <= 1'd0;
		vns_new_master_wdata_ready4 <= 1'd0;
		vns_new_master_wdata_ready5 <= 1'd0;
		vns_new_master_wdata_ready6 <= 1'd0;
		vns_new_master_wdata_ready7 <= 1'd0;
		vns_new_master_wdata_ready8 <= 1'd0;
		vns_new_master_rdata_valid0 <= 1'd0;
		vns_new_master_rdata_valid1 <= 1'd0;
		vns_new_master_rdata_valid2 <= 1'd0;
		vns_new_master_rdata_valid3 <= 1'd0;
		vns_new_master_rdata_valid4 <= 1'd0;
		vns_new_master_rdata_valid5 <= 1'd0;
		vns_new_master_rdata_valid6 <= 1'd0;
		vns_new_master_rdata_valid7 <= 1'd0;
		vns_new_master_rdata_valid8 <= 1'd0;
		vns_new_master_rdata_valid9 <= 1'd0;
		vns_new_master_rdata_valid10 <= 1'd0;
		vns_new_master_rdata_valid11 <= 1'd0;
		vns_new_master_rdata_valid12 <= 1'd0;
		vns_new_master_rdata_valid13 <= 1'd0;
		vns_new_master_rdata_valid14 <= 1'd0;
		vns_new_master_rdata_valid15 <= 1'd0;
		vns_new_master_rdata_valid16 <= 1'd0;
		vns_new_master_rdata_valid17 <= 1'd0;
		vns_new_master_rdata_valid18 <= 1'd0;
		vns_new_master_rdata_valid19 <= 1'd0;
		vns_new_master_rdata_valid20 <= 1'd0;
		vns_fullmemorywe_state <= 3'd0;
		vns_litedramwishbonebridge_state <= 2'd0;
		vns_liteethmacsramwriter_state <= 2'd0;
		vns_liteethmacsramreader_state <= 2'd0;
		vns_edid_state <= 4'd0;
		vns_dma_state <= 2'd0;
		vns_videosoc_grant <= 2'd0;
		vns_videosoc_slave_sel_r <= 6'd0;
		vns_videosoc_interface0_bank_bus_dat_r <= 8'd0;
		vns_videosoc_interface1_bank_bus_dat_r <= 8'd0;
		vns_videosoc_interface2_bank_bus_dat_r <= 8'd0;
		vns_videosoc_sel_r <= 1'd0;
		vns_videosoc_interface3_bank_bus_dat_r <= 8'd0;
		vns_videosoc_interface4_bank_bus_dat_r <= 8'd0;
		vns_videosoc_interface5_bank_bus_dat_r <= 8'd0;
		vns_videosoc_csrbank5_core_initiator_hres_backstore <= 4'd0;
		vns_videosoc_csrbank5_core_initiator_hsync_start_backstore <= 4'd0;
		vns_videosoc_csrbank5_core_initiator_hsync_end_backstore <= 4'd0;
		vns_videosoc_csrbank5_core_initiator_hscan_backstore <= 4'd0;
		vns_videosoc_csrbank5_core_initiator_vres_backstore <= 4'd0;
		vns_videosoc_csrbank5_core_initiator_vsync_start_backstore <= 4'd0;
		vns_videosoc_csrbank5_core_initiator_vsync_end_backstore <= 4'd0;
		vns_videosoc_csrbank5_core_initiator_vscan_backstore <= 4'd0;
		vns_videosoc_csrbank5_core_initiator_base_backstore <= 24'd0;
		vns_videosoc_csrbank5_core_initiator_length_backstore <= 24'd0;
		vns_videosoc_interface6_bank_bus_dat_r <= 8'd0;
		vns_videosoc_interface7_bank_bus_dat_r <= 8'd0;
		vns_videosoc_interface8_bank_bus_dat_r <= 8'd0;
		vns_videosoc_interface9_bank_bus_dat_r <= 8'd0;
		vns_videosoc_interface10_bank_bus_dat_r <= 8'd0;
		vns_videosoc_interface11_bank_bus_dat_r <= 8'd0;
		vns_videosoc_interface12_bank_bus_dat_r <= 8'd0;
	end
	vns_xilinxmultiregimpl0_regs0 <= serial_rx;
	vns_xilinxmultiregimpl0_regs1 <= vns_xilinxmultiregimpl0_regs0;
	vns_xilinxmultiregimpl1_regs0 <= soc_ethphy_data_r;
	vns_xilinxmultiregimpl1_regs1 <= vns_xilinxmultiregimpl1_regs0;
	vns_xilinxmultiregimpl3_regs0 <= soc_ethmac_tx_cdc_graycounter1_q;
	vns_xilinxmultiregimpl3_regs1 <= vns_xilinxmultiregimpl3_regs0;
	vns_xilinxmultiregimpl4_regs0 <= soc_ethmac_rx_cdc_graycounter0_q;
	vns_xilinxmultiregimpl4_regs1 <= vns_xilinxmultiregimpl4_regs0;
	vns_xilinxmultiregimpl6_regs0 <= hdmi_in_scl;
	vns_xilinxmultiregimpl6_regs1 <= vns_xilinxmultiregimpl6_regs0;
	vns_xilinxmultiregimpl7_regs0 <= soc_edid_sda_i_async;
	vns_xilinxmultiregimpl7_regs1 <= vns_xilinxmultiregimpl7_regs0;
	vns_xilinxmultiregimpl8_regs0 <= soc_mmcm_locked;
	vns_xilinxmultiregimpl8_regs1 <= vns_xilinxmultiregimpl8_regs0;
	vns_xilinxmultiregimpl14_regs0 <= {soc_s7datacapture0_too_early, soc_s7datacapture0_too_late};
	vns_xilinxmultiregimpl14_regs1 <= vns_xilinxmultiregimpl14_regs0;
	vns_xilinxmultiregimpl16_regs0 <= soc_charsync0_synced;
	vns_xilinxmultiregimpl16_regs1 <= vns_xilinxmultiregimpl16_regs0;
	vns_xilinxmultiregimpl17_regs0 <= soc_charsync0_word_sel;
	vns_xilinxmultiregimpl17_regs1 <= vns_xilinxmultiregimpl17_regs0;
	vns_xilinxmultiregimpl18_regs0 <= soc_wer0_toggle_i;
	vns_xilinxmultiregimpl18_regs1 <= vns_xilinxmultiregimpl18_regs0;
	vns_xilinxmultiregimpl24_regs0 <= {soc_s7datacapture1_too_early, soc_s7datacapture1_too_late};
	vns_xilinxmultiregimpl24_regs1 <= vns_xilinxmultiregimpl24_regs0;
	vns_xilinxmultiregimpl26_regs0 <= soc_charsync1_synced;
	vns_xilinxmultiregimpl26_regs1 <= vns_xilinxmultiregimpl26_regs0;
	vns_xilinxmultiregimpl27_regs0 <= soc_charsync1_word_sel;
	vns_xilinxmultiregimpl27_regs1 <= vns_xilinxmultiregimpl27_regs0;
	vns_xilinxmultiregimpl28_regs0 <= soc_wer1_toggle_i;
	vns_xilinxmultiregimpl28_regs1 <= vns_xilinxmultiregimpl28_regs0;
	vns_xilinxmultiregimpl34_regs0 <= {soc_s7datacapture2_too_early, soc_s7datacapture2_too_late};
	vns_xilinxmultiregimpl34_regs1 <= vns_xilinxmultiregimpl34_regs0;
	vns_xilinxmultiregimpl36_regs0 <= soc_charsync2_synced;
	vns_xilinxmultiregimpl36_regs1 <= vns_xilinxmultiregimpl36_regs0;
	vns_xilinxmultiregimpl37_regs0 <= soc_charsync2_word_sel;
	vns_xilinxmultiregimpl37_regs1 <= vns_xilinxmultiregimpl37_regs0;
	vns_xilinxmultiregimpl38_regs0 <= soc_wer2_toggle_i;
	vns_xilinxmultiregimpl38_regs1 <= vns_xilinxmultiregimpl38_regs0;
	vns_xilinxmultiregimpl39_regs0 <= soc_chansync_chan_synced;
	vns_xilinxmultiregimpl39_regs1 <= vns_xilinxmultiregimpl39_regs0;
	vns_xilinxmultiregimpl40_regs0 <= soc_resdetection_hcounter_st;
	vns_xilinxmultiregimpl40_regs1 <= vns_xilinxmultiregimpl40_regs0;
	vns_xilinxmultiregimpl41_regs0 <= soc_resdetection_vcounter_st;
	vns_xilinxmultiregimpl41_regs1 <= vns_xilinxmultiregimpl41_regs0;
	vns_xilinxmultiregimpl42_regs0 <= soc_frame_fifo_graycounter0_q;
	vns_xilinxmultiregimpl42_regs1 <= vns_xilinxmultiregimpl42_regs0;
	vns_xilinxmultiregimpl44_regs0 <= soc_frame_pix_overflow;
	vns_xilinxmultiregimpl44_regs1 <= vns_xilinxmultiregimpl44_regs0;
	vns_xilinxmultiregimpl46_regs0 <= soc_frame_overflow_reset_ack_toggle_i;
	vns_xilinxmultiregimpl46_regs1 <= vns_xilinxmultiregimpl46_regs0;
	vns_xilinxmultiregimpl47_regs0 <= soc_hdmi_in0_freq_q;
	vns_xilinxmultiregimpl47_regs1 <= vns_xilinxmultiregimpl47_regs0;
	vns_xilinxmultiregimpl48_regs0 <= soc_hdmi_out0_dram_port_cmd_fifo_graycounter0_q;
	vns_xilinxmultiregimpl48_regs1 <= vns_xilinxmultiregimpl48_regs0;
	vns_xilinxmultiregimpl51_regs0 <= soc_hdmi_out0_dram_port_rdata_fifo_graycounter1_q;
	vns_xilinxmultiregimpl51_regs1 <= vns_xilinxmultiregimpl51_regs0;
	vns_xilinxmultiregimpl53_regs0 <= soc_hdmi_out0_core_initiator_cdc_graycounter1_q;
	vns_xilinxmultiregimpl53_regs1 <= vns_xilinxmultiregimpl53_regs0;
	vns_xilinxmultiregimpl54_regs0 <= soc_hdmi_out0_core_underflow_enable_storage;
	vns_xilinxmultiregimpl54_regs1 <= vns_xilinxmultiregimpl54_regs0;
end

lm32_cpu #(
	.eba_reset(32'h00000000)
) lm32_cpu (
	.D_ACK_I(soc_videosoc_videosoc_dbus_ack),
	.D_DAT_I(soc_videosoc_videosoc_dbus_dat_r),
	.D_ERR_I(soc_videosoc_videosoc_dbus_err),
	.D_RTY_I(1'd0),
	.I_ACK_I(soc_videosoc_videosoc_ibus_ack),
	.I_DAT_I(soc_videosoc_videosoc_ibus_dat_r),
	.I_ERR_I(soc_videosoc_videosoc_ibus_err),
	.I_RTY_I(1'd0),
	.clk_i(sys_clk),
	.interrupt(soc_videosoc_videosoc_interrupt),
	.rst_i(sys_rst),
	.D_ADR_O(soc_videosoc_videosoc_d_adr_o),
	.D_BTE_O(soc_videosoc_videosoc_dbus_bte),
	.D_CTI_O(soc_videosoc_videosoc_dbus_cti),
	.D_CYC_O(soc_videosoc_videosoc_dbus_cyc),
	.D_DAT_O(soc_videosoc_videosoc_dbus_dat_w),
	.D_SEL_O(soc_videosoc_videosoc_dbus_sel),
	.D_STB_O(soc_videosoc_videosoc_dbus_stb),
	.D_WE_O(soc_videosoc_videosoc_dbus_we),
	.I_ADR_O(soc_videosoc_videosoc_i_adr_o),
	.I_BTE_O(soc_videosoc_videosoc_ibus_bte),
	.I_CTI_O(soc_videosoc_videosoc_ibus_cti),
	.I_CYC_O(soc_videosoc_videosoc_ibus_cyc),
	.I_DAT_O(soc_videosoc_videosoc_ibus_dat_w),
	.I_SEL_O(soc_videosoc_videosoc_ibus_sel),
	.I_STB_O(soc_videosoc_videosoc_ibus_stb),
	.I_WE_O(soc_videosoc_videosoc_ibus_we)
);

reg [31:0] mem[0:8191];
reg [31:0] memdat;
always @(posedge sys_clk) begin
	memdat <= mem[soc_videosoc_videosoc_rom_adr];
end

assign soc_videosoc_videosoc_rom_dat_r = memdat;

initial begin
	$readmemh("mem.init", mem);
end

reg [31:0] mem_1[0:8191];
reg [12:0] memadr;
always @(posedge sys_clk) begin
	if (soc_videosoc_videosoc_sram_we[0])
		mem_1[soc_videosoc_videosoc_sram_adr][7:0] <= soc_videosoc_videosoc_sram_dat_w[7:0];
	if (soc_videosoc_videosoc_sram_we[1])
		mem_1[soc_videosoc_videosoc_sram_adr][15:8] <= soc_videosoc_videosoc_sram_dat_w[15:8];
	if (soc_videosoc_videosoc_sram_we[2])
		mem_1[soc_videosoc_videosoc_sram_adr][23:16] <= soc_videosoc_videosoc_sram_dat_w[23:16];
	if (soc_videosoc_videosoc_sram_we[3])
		mem_1[soc_videosoc_videosoc_sram_adr][31:24] <= soc_videosoc_videosoc_sram_dat_w[31:24];
	memadr <= soc_videosoc_videosoc_sram_adr;
end

assign soc_videosoc_videosoc_sram_dat_r = mem_1[memadr];

PLLE2_BASE #(
	.CLKFBOUT_MULT(5'd16),
	.CLKIN1_PERIOD(10.0),
	.CLKOUT0_DIVIDE(5'd16),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(3'd4),
	.CLKOUT1_PHASE(0.0),
	.CLKOUT2_DIVIDE(3'd4),
	.CLKOUT2_PHASE(90.0),
	.CLKOUT3_DIVIDE(4'd8),
	.CLKOUT3_PHASE(0.0),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER1(0.01),
	.STARTUP_WAIT("FALSE")
) PLLE2_BASE (
	.CLKFBIN(soc_videosoc_pll_fb),
	.CLKIN1(clk100),
	.CLKFBOUT(soc_videosoc_pll_fb),
	.CLKOUT0(soc_videosoc_pll_sys),
	.CLKOUT1(soc_videosoc_pll_sys4x),
	.CLKOUT2(soc_videosoc_pll_sys4x_dqs),
	.CLKOUT3(soc_videosoc_pll_clk200),
	.LOCKED(soc_videosoc_pll_locked)
);

BUFG BUFG(
	.I(soc_videosoc_pll_sys),
	.O(sys_clk)
);

BUFG BUFG_1(
	.I(soc_videosoc_pll_sys4x),
	.O(sys4x_clk)
);

BUFG BUFG_2(
	.I(soc_videosoc_pll_sys4x_dqs),
	.O(sys4x_dqs_clk)
);

BUFG BUFG_3(
	.I(soc_videosoc_pll_clk200),
	.O(clk200_clk)
);

BUFG BUFG_4(
	.I(clk100),
	.O(clk100_clk)
);

IDELAYCTRL IDELAYCTRL(
	.REFCLK(clk200_clk),
	.RST(soc_videosoc_ic_reset)
);

reg [9:0] storage[0:15];
reg [3:0] memadr_1;
always @(posedge sys_clk) begin
	if (soc_videosoc_uart_tx_fifo_wrport_we)
		storage[soc_videosoc_uart_tx_fifo_wrport_adr] <= soc_videosoc_uart_tx_fifo_wrport_dat_w;
	memadr_1 <= soc_videosoc_uart_tx_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign soc_videosoc_uart_tx_fifo_wrport_dat_r = storage[memadr_1];
assign soc_videosoc_uart_tx_fifo_rdport_dat_r = storage[soc_videosoc_uart_tx_fifo_rdport_adr];

reg [9:0] storage_1[0:15];
reg [3:0] memadr_2;
always @(posedge sys_clk) begin
	if (soc_videosoc_uart_rx_fifo_wrport_we)
		storage_1[soc_videosoc_uart_rx_fifo_wrport_adr] <= soc_videosoc_uart_rx_fifo_wrport_dat_w;
	memadr_2 <= soc_videosoc_uart_rx_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign soc_videosoc_uart_rx_fifo_wrport_dat_r = storage_1[memadr_2];
assign soc_videosoc_uart_rx_fifo_rdport_dat_r = storage_1[soc_videosoc_uart_rx_fifo_rdport_adr];

DNA_PORT DNA_PORT(
	.CLK(soc_videosoc_info_dna_cnt[0]),
	.DIN(soc_videosoc_info_dna_status[56]),
	.READ((soc_videosoc_info_dna_cnt < 2'd2)),
	.SHIFT(1'd1),
	.DOUT(soc_videosoc_info_dna_do)
);

XADC #(
	.INIT_40(16'd36864),
	.INIT_41(14'd12016),
	.INIT_42(11'd1024),
	.INIT_48(15'd18177),
	.INIT_49(4'd15),
	.INIT_4A(15'd18176),
	.INIT_4B(1'd0),
	.INIT_4C(1'd0),
	.INIT_4D(1'd0),
	.INIT_4E(1'd0),
	.INIT_4F(1'd0),
	.INIT_50(16'd46573),
	.INIT_51(15'd22937),
	.INIT_52(16'd41287),
	.INIT_53(16'd56797),
	.INIT_54(16'd43322),
	.INIT_55(15'd20753),
	.INIT_56(16'd37355),
	.INIT_57(16'd44622),
	.INIT_58(15'd22937),
	.INIT_5C(15'd20753)
) XADC (
	.CONVST(1'd0),
	.CONVSTCLK(1'd0),
	.DADDR(soc_videosoc_info_channel),
	.DCLK(sys_clk),
	.DEN(soc_videosoc_info_eoc),
	.DI(1'd0),
	.DWE(1'd0),
	.RESET(sys_rst),
	.VAUXN(1'd0),
	.VAUXP(1'd1),
	.VN(1'd0),
	.VP(1'd1),
	.ALM(soc_videosoc_info_alarm),
	.BUSY(soc_videosoc_info_busy),
	.CHANNEL(soc_videosoc_info_channel),
	.DO(soc_videosoc_info_data),
	.DRDY(soc_videosoc_info_drdy),
	.EOC(soc_videosoc_info_eoc),
	.EOS(soc_videosoc_info_eos),
	.OT(soc_videosoc_info_ot)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(1'd0),
	.D2(1'd1),
	.D3(1'd0),
	.D4(1'd1),
	.D5(1'd0),
	.D6(1'd1),
	.D7(1'd0),
	.D8(1'd1),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(soc_videosoc_ddrphy_sd_clk_se)
);

OBUFDS OBUFDS(
	.I(soc_videosoc_ddrphy_sd_clk_se),
	.O(ddram_clk_p),
	.OB(ddram_clk_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_1 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_address[0]),
	.D2(soc_videosoc_ddrphy_dfi_p0_address[0]),
	.D3(soc_videosoc_ddrphy_dfi_p1_address[0]),
	.D4(soc_videosoc_ddrphy_dfi_p1_address[0]),
	.D5(soc_videosoc_ddrphy_dfi_p2_address[0]),
	.D6(soc_videosoc_ddrphy_dfi_p2_address[0]),
	.D7(soc_videosoc_ddrphy_dfi_p3_address[0]),
	.D8(soc_videosoc_ddrphy_dfi_p3_address[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_address[1]),
	.D2(soc_videosoc_ddrphy_dfi_p0_address[1]),
	.D3(soc_videosoc_ddrphy_dfi_p1_address[1]),
	.D4(soc_videosoc_ddrphy_dfi_p1_address[1]),
	.D5(soc_videosoc_ddrphy_dfi_p2_address[1]),
	.D6(soc_videosoc_ddrphy_dfi_p2_address[1]),
	.D7(soc_videosoc_ddrphy_dfi_p3_address[1]),
	.D8(soc_videosoc_ddrphy_dfi_p3_address[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_3 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_address[2]),
	.D2(soc_videosoc_ddrphy_dfi_p0_address[2]),
	.D3(soc_videosoc_ddrphy_dfi_p1_address[2]),
	.D4(soc_videosoc_ddrphy_dfi_p1_address[2]),
	.D5(soc_videosoc_ddrphy_dfi_p2_address[2]),
	.D6(soc_videosoc_ddrphy_dfi_p2_address[2]),
	.D7(soc_videosoc_ddrphy_dfi_p3_address[2]),
	.D8(soc_videosoc_ddrphy_dfi_p3_address[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_4 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_address[3]),
	.D2(soc_videosoc_ddrphy_dfi_p0_address[3]),
	.D3(soc_videosoc_ddrphy_dfi_p1_address[3]),
	.D4(soc_videosoc_ddrphy_dfi_p1_address[3]),
	.D5(soc_videosoc_ddrphy_dfi_p2_address[3]),
	.D6(soc_videosoc_ddrphy_dfi_p2_address[3]),
	.D7(soc_videosoc_ddrphy_dfi_p3_address[3]),
	.D8(soc_videosoc_ddrphy_dfi_p3_address[3]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[3])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_5 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_address[4]),
	.D2(soc_videosoc_ddrphy_dfi_p0_address[4]),
	.D3(soc_videosoc_ddrphy_dfi_p1_address[4]),
	.D4(soc_videosoc_ddrphy_dfi_p1_address[4]),
	.D5(soc_videosoc_ddrphy_dfi_p2_address[4]),
	.D6(soc_videosoc_ddrphy_dfi_p2_address[4]),
	.D7(soc_videosoc_ddrphy_dfi_p3_address[4]),
	.D8(soc_videosoc_ddrphy_dfi_p3_address[4]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[4])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_6 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_address[5]),
	.D2(soc_videosoc_ddrphy_dfi_p0_address[5]),
	.D3(soc_videosoc_ddrphy_dfi_p1_address[5]),
	.D4(soc_videosoc_ddrphy_dfi_p1_address[5]),
	.D5(soc_videosoc_ddrphy_dfi_p2_address[5]),
	.D6(soc_videosoc_ddrphy_dfi_p2_address[5]),
	.D7(soc_videosoc_ddrphy_dfi_p3_address[5]),
	.D8(soc_videosoc_ddrphy_dfi_p3_address[5]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[5])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_7 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_address[6]),
	.D2(soc_videosoc_ddrphy_dfi_p0_address[6]),
	.D3(soc_videosoc_ddrphy_dfi_p1_address[6]),
	.D4(soc_videosoc_ddrphy_dfi_p1_address[6]),
	.D5(soc_videosoc_ddrphy_dfi_p2_address[6]),
	.D6(soc_videosoc_ddrphy_dfi_p2_address[6]),
	.D7(soc_videosoc_ddrphy_dfi_p3_address[6]),
	.D8(soc_videosoc_ddrphy_dfi_p3_address[6]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[6])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_8 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_address[7]),
	.D2(soc_videosoc_ddrphy_dfi_p0_address[7]),
	.D3(soc_videosoc_ddrphy_dfi_p1_address[7]),
	.D4(soc_videosoc_ddrphy_dfi_p1_address[7]),
	.D5(soc_videosoc_ddrphy_dfi_p2_address[7]),
	.D6(soc_videosoc_ddrphy_dfi_p2_address[7]),
	.D7(soc_videosoc_ddrphy_dfi_p3_address[7]),
	.D8(soc_videosoc_ddrphy_dfi_p3_address[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[7])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_9 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_address[8]),
	.D2(soc_videosoc_ddrphy_dfi_p0_address[8]),
	.D3(soc_videosoc_ddrphy_dfi_p1_address[8]),
	.D4(soc_videosoc_ddrphy_dfi_p1_address[8]),
	.D5(soc_videosoc_ddrphy_dfi_p2_address[8]),
	.D6(soc_videosoc_ddrphy_dfi_p2_address[8]),
	.D7(soc_videosoc_ddrphy_dfi_p3_address[8]),
	.D8(soc_videosoc_ddrphy_dfi_p3_address[8]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[8])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_10 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_address[9]),
	.D2(soc_videosoc_ddrphy_dfi_p0_address[9]),
	.D3(soc_videosoc_ddrphy_dfi_p1_address[9]),
	.D4(soc_videosoc_ddrphy_dfi_p1_address[9]),
	.D5(soc_videosoc_ddrphy_dfi_p2_address[9]),
	.D6(soc_videosoc_ddrphy_dfi_p2_address[9]),
	.D7(soc_videosoc_ddrphy_dfi_p3_address[9]),
	.D8(soc_videosoc_ddrphy_dfi_p3_address[9]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[9])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_11 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_address[10]),
	.D2(soc_videosoc_ddrphy_dfi_p0_address[10]),
	.D3(soc_videosoc_ddrphy_dfi_p1_address[10]),
	.D4(soc_videosoc_ddrphy_dfi_p1_address[10]),
	.D5(soc_videosoc_ddrphy_dfi_p2_address[10]),
	.D6(soc_videosoc_ddrphy_dfi_p2_address[10]),
	.D7(soc_videosoc_ddrphy_dfi_p3_address[10]),
	.D8(soc_videosoc_ddrphy_dfi_p3_address[10]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[10])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_12 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_address[11]),
	.D2(soc_videosoc_ddrphy_dfi_p0_address[11]),
	.D3(soc_videosoc_ddrphy_dfi_p1_address[11]),
	.D4(soc_videosoc_ddrphy_dfi_p1_address[11]),
	.D5(soc_videosoc_ddrphy_dfi_p2_address[11]),
	.D6(soc_videosoc_ddrphy_dfi_p2_address[11]),
	.D7(soc_videosoc_ddrphy_dfi_p3_address[11]),
	.D8(soc_videosoc_ddrphy_dfi_p3_address[11]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[11])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_13 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_address[12]),
	.D2(soc_videosoc_ddrphy_dfi_p0_address[12]),
	.D3(soc_videosoc_ddrphy_dfi_p1_address[12]),
	.D4(soc_videosoc_ddrphy_dfi_p1_address[12]),
	.D5(soc_videosoc_ddrphy_dfi_p2_address[12]),
	.D6(soc_videosoc_ddrphy_dfi_p2_address[12]),
	.D7(soc_videosoc_ddrphy_dfi_p3_address[12]),
	.D8(soc_videosoc_ddrphy_dfi_p3_address[12]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[12])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_14 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_address[13]),
	.D2(soc_videosoc_ddrphy_dfi_p0_address[13]),
	.D3(soc_videosoc_ddrphy_dfi_p1_address[13]),
	.D4(soc_videosoc_ddrphy_dfi_p1_address[13]),
	.D5(soc_videosoc_ddrphy_dfi_p2_address[13]),
	.D6(soc_videosoc_ddrphy_dfi_p2_address[13]),
	.D7(soc_videosoc_ddrphy_dfi_p3_address[13]),
	.D8(soc_videosoc_ddrphy_dfi_p3_address[13]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[13])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_15 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_address[14]),
	.D2(soc_videosoc_ddrphy_dfi_p0_address[14]),
	.D3(soc_videosoc_ddrphy_dfi_p1_address[14]),
	.D4(soc_videosoc_ddrphy_dfi_p1_address[14]),
	.D5(soc_videosoc_ddrphy_dfi_p2_address[14]),
	.D6(soc_videosoc_ddrphy_dfi_p2_address[14]),
	.D7(soc_videosoc_ddrphy_dfi_p3_address[14]),
	.D8(soc_videosoc_ddrphy_dfi_p3_address[14]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a[14])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_16 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_bank[0]),
	.D2(soc_videosoc_ddrphy_dfi_p0_bank[0]),
	.D3(soc_videosoc_ddrphy_dfi_p1_bank[0]),
	.D4(soc_videosoc_ddrphy_dfi_p1_bank[0]),
	.D5(soc_videosoc_ddrphy_dfi_p2_bank[0]),
	.D6(soc_videosoc_ddrphy_dfi_p2_bank[0]),
	.D7(soc_videosoc_ddrphy_dfi_p3_bank[0]),
	.D8(soc_videosoc_ddrphy_dfi_p3_bank[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_17 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_bank[1]),
	.D2(soc_videosoc_ddrphy_dfi_p0_bank[1]),
	.D3(soc_videosoc_ddrphy_dfi_p1_bank[1]),
	.D4(soc_videosoc_ddrphy_dfi_p1_bank[1]),
	.D5(soc_videosoc_ddrphy_dfi_p2_bank[1]),
	.D6(soc_videosoc_ddrphy_dfi_p2_bank[1]),
	.D7(soc_videosoc_ddrphy_dfi_p3_bank[1]),
	.D8(soc_videosoc_ddrphy_dfi_p3_bank[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_18 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_bank[2]),
	.D2(soc_videosoc_ddrphy_dfi_p0_bank[2]),
	.D3(soc_videosoc_ddrphy_dfi_p1_bank[2]),
	.D4(soc_videosoc_ddrphy_dfi_p1_bank[2]),
	.D5(soc_videosoc_ddrphy_dfi_p2_bank[2]),
	.D6(soc_videosoc_ddrphy_dfi_p2_bank[2]),
	.D7(soc_videosoc_ddrphy_dfi_p3_bank[2]),
	.D8(soc_videosoc_ddrphy_dfi_p3_bank[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba[2])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_19 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_ras_n),
	.D2(soc_videosoc_ddrphy_dfi_p0_ras_n),
	.D3(soc_videosoc_ddrphy_dfi_p1_ras_n),
	.D4(soc_videosoc_ddrphy_dfi_p1_ras_n),
	.D5(soc_videosoc_ddrphy_dfi_p2_ras_n),
	.D6(soc_videosoc_ddrphy_dfi_p2_ras_n),
	.D7(soc_videosoc_ddrphy_dfi_p3_ras_n),
	.D8(soc_videosoc_ddrphy_dfi_p3_ras_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ras_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_20 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_cas_n),
	.D2(soc_videosoc_ddrphy_dfi_p0_cas_n),
	.D3(soc_videosoc_ddrphy_dfi_p1_cas_n),
	.D4(soc_videosoc_ddrphy_dfi_p1_cas_n),
	.D5(soc_videosoc_ddrphy_dfi_p2_cas_n),
	.D6(soc_videosoc_ddrphy_dfi_p2_cas_n),
	.D7(soc_videosoc_ddrphy_dfi_p3_cas_n),
	.D8(soc_videosoc_ddrphy_dfi_p3_cas_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cas_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_21 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_we_n),
	.D2(soc_videosoc_ddrphy_dfi_p0_we_n),
	.D3(soc_videosoc_ddrphy_dfi_p1_we_n),
	.D4(soc_videosoc_ddrphy_dfi_p1_we_n),
	.D5(soc_videosoc_ddrphy_dfi_p2_we_n),
	.D6(soc_videosoc_ddrphy_dfi_p2_we_n),
	.D7(soc_videosoc_ddrphy_dfi_p3_we_n),
	.D8(soc_videosoc_ddrphy_dfi_p3_we_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_we_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_22 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_cke),
	.D2(soc_videosoc_ddrphy_dfi_p0_cke),
	.D3(soc_videosoc_ddrphy_dfi_p1_cke),
	.D4(soc_videosoc_ddrphy_dfi_p1_cke),
	.D5(soc_videosoc_ddrphy_dfi_p2_cke),
	.D6(soc_videosoc_ddrphy_dfi_p2_cke),
	.D7(soc_videosoc_ddrphy_dfi_p3_cke),
	.D8(soc_videosoc_ddrphy_dfi_p3_cke),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cke)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_23 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_odt),
	.D2(soc_videosoc_ddrphy_dfi_p0_odt),
	.D3(soc_videosoc_ddrphy_dfi_p1_odt),
	.D4(soc_videosoc_ddrphy_dfi_p1_odt),
	.D5(soc_videosoc_ddrphy_dfi_p2_odt),
	.D6(soc_videosoc_ddrphy_dfi_p2_odt),
	.D7(soc_videosoc_ddrphy_dfi_p3_odt),
	.D8(soc_videosoc_ddrphy_dfi_p3_odt),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_odt)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_24 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_reset_n),
	.D2(soc_videosoc_ddrphy_dfi_p0_reset_n),
	.D3(soc_videosoc_ddrphy_dfi_p1_reset_n),
	.D4(soc_videosoc_ddrphy_dfi_p1_reset_n),
	.D5(soc_videosoc_ddrphy_dfi_p2_reset_n),
	.D6(soc_videosoc_ddrphy_dfi_p2_reset_n),
	.D7(soc_videosoc_ddrphy_dfi_p3_reset_n),
	.D8(soc_videosoc_ddrphy_dfi_p3_reset_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_reset_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_25 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata_mask[0]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata_mask[2]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata_mask[0]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata_mask[2]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata_mask[0]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata_mask[2]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata_mask[0]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata_mask[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_26 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dqs_serdes_pattern[0]),
	.D2(soc_videosoc_ddrphy_dqs_serdes_pattern[1]),
	.D3(soc_videosoc_ddrphy_dqs_serdes_pattern[2]),
	.D4(soc_videosoc_ddrphy_dqs_serdes_pattern[3]),
	.D5(soc_videosoc_ddrphy_dqs_serdes_pattern[4]),
	.D6(soc_videosoc_ddrphy_dqs_serdes_pattern[5]),
	.D7(soc_videosoc_ddrphy_dqs_serdes_pattern[6]),
	.D8(soc_videosoc_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dqs0),
	.TQ(soc_videosoc_ddrphy_dqs_t0)
);

OBUFTDS OBUFTDS(
	.I(soc_videosoc_ddrphy_dqs0),
	.T(soc_videosoc_ddrphy_dqs_t0),
	.O(ddram_dqs_p[0]),
	.OB(ddram_dqs_n[0])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_27 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata_mask[1]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata_mask[3]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata_mask[1]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata_mask[3]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata_mask[1]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata_mask[3]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata_mask[1]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata_mask[3]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_28 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dqs_serdes_pattern[0]),
	.D2(soc_videosoc_ddrphy_dqs_serdes_pattern[1]),
	.D3(soc_videosoc_ddrphy_dqs_serdes_pattern[2]),
	.D4(soc_videosoc_ddrphy_dqs_serdes_pattern[3]),
	.D5(soc_videosoc_ddrphy_dqs_serdes_pattern[4]),
	.D6(soc_videosoc_ddrphy_dqs_serdes_pattern[5]),
	.D7(soc_videosoc_ddrphy_dqs_serdes_pattern[6]),
	.D8(soc_videosoc_ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dqs1),
	.TQ(soc_videosoc_ddrphy_dqs_t1)
);

OBUFTDS OBUFTDS_1(
	.I(soc_videosoc_ddrphy_dqs1),
	.T(soc_videosoc_ddrphy_dqs_t1),
	.O(ddram_dqs_p[1]),
	.OB(ddram_dqs_n[1])
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_29 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[0]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[16]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[0]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[16]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[0]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[16]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[0]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[16]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o0),
	.TQ(soc_videosoc_ddrphy_dq_t0)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2 (
	.BITSLIP((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed0),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[16]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[0]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[16]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[0]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[16]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[0]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[16]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay0),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed0)
);

IOBUF IOBUF(
	.I(soc_videosoc_ddrphy_dq_o0),
	.T(soc_videosoc_ddrphy_dq_t0),
	.IO(ddram_dq[0]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay0)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_30 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[1]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[17]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[1]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[17]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[1]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[17]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[1]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[17]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o1),
	.TQ(soc_videosoc_ddrphy_dq_t1)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_1 (
	.BITSLIP((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed1),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[17]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[1]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[17]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[1]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[17]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[1]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[17]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[1])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_1 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay1),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed1)
);

IOBUF IOBUF_1(
	.I(soc_videosoc_ddrphy_dq_o1),
	.T(soc_videosoc_ddrphy_dq_t1),
	.IO(ddram_dq[1]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay1)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_31 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[2]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[18]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[2]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[18]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[2]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[18]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[2]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[18]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o2),
	.TQ(soc_videosoc_ddrphy_dq_t2)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_2 (
	.BITSLIP((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed2),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[18]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[2]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[18]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[2]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[18]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[2]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[18]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[2])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_2 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay2),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed2)
);

IOBUF IOBUF_2(
	.I(soc_videosoc_ddrphy_dq_o2),
	.T(soc_videosoc_ddrphy_dq_t2),
	.IO(ddram_dq[2]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay2)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_32 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[3]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[19]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[3]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[19]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[3]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[19]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[3]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[19]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o3),
	.TQ(soc_videosoc_ddrphy_dq_t3)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_3 (
	.BITSLIP((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed3),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[19]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[3]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[19]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[3]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[19]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[3]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[19]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[3])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_3 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay3),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed3)
);

IOBUF IOBUF_3(
	.I(soc_videosoc_ddrphy_dq_o3),
	.T(soc_videosoc_ddrphy_dq_t3),
	.IO(ddram_dq[3]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay3)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_33 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[4]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[20]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[4]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[20]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[4]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[20]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[4]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[20]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o4),
	.TQ(soc_videosoc_ddrphy_dq_t4)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_4 (
	.BITSLIP((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed4),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[20]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[4]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[20]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[4]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[20]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[4]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[20]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[4])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_4 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay4),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed4)
);

IOBUF IOBUF_4(
	.I(soc_videosoc_ddrphy_dq_o4),
	.T(soc_videosoc_ddrphy_dq_t4),
	.IO(ddram_dq[4]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay4)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_34 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[5]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[21]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[5]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[21]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[5]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[21]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[5]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[21]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o5),
	.TQ(soc_videosoc_ddrphy_dq_t5)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_5 (
	.BITSLIP((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed5),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[21]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[5]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[21]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[5]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[21]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[5]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[21]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[5])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_5 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay5),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed5)
);

IOBUF IOBUF_5(
	.I(soc_videosoc_ddrphy_dq_o5),
	.T(soc_videosoc_ddrphy_dq_t5),
	.IO(ddram_dq[5]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay5)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_35 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[6]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[22]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[6]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[22]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[6]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[22]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[6]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[22]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o6),
	.TQ(soc_videosoc_ddrphy_dq_t6)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_6 (
	.BITSLIP((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed6),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[22]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[6]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[22]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[6]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[22]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[6]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[22]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[6])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_6 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay6),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed6)
);

IOBUF IOBUF_6(
	.I(soc_videosoc_ddrphy_dq_o6),
	.T(soc_videosoc_ddrphy_dq_t6),
	.IO(ddram_dq[6]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay6)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_36 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[7]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[23]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[7]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[23]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[7]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[23]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[7]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[23]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o7),
	.TQ(soc_videosoc_ddrphy_dq_t7)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_7 (
	.BITSLIP((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed7),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[23]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[7]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[23]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[7]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[23]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[7]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[23]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[7])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_7 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay7),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[0] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed7)
);

IOBUF IOBUF_7(
	.I(soc_videosoc_ddrphy_dq_o7),
	.T(soc_videosoc_ddrphy_dq_t7),
	.IO(ddram_dq[7]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay7)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_37 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[8]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[24]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[8]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[24]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[8]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[24]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[8]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[24]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o8),
	.TQ(soc_videosoc_ddrphy_dq_t8)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_8 (
	.BITSLIP((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed8),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[24]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[8]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[24]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[8]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[24]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[8]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[24]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[8])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_8 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay8),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed8)
);

IOBUF IOBUF_8(
	.I(soc_videosoc_ddrphy_dq_o8),
	.T(soc_videosoc_ddrphy_dq_t8),
	.IO(ddram_dq[8]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay8)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_38 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[9]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[25]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[9]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[25]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[9]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[25]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[9]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[25]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o9),
	.TQ(soc_videosoc_ddrphy_dq_t9)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_9 (
	.BITSLIP((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed9),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[25]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[9]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[25]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[9]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[25]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[9]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[25]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[9])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_9 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay9),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed9)
);

IOBUF IOBUF_9(
	.I(soc_videosoc_ddrphy_dq_o9),
	.T(soc_videosoc_ddrphy_dq_t9),
	.IO(ddram_dq[9]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay9)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_39 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[10]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[26]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[10]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[26]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[10]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[26]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[10]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[26]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o10),
	.TQ(soc_videosoc_ddrphy_dq_t10)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_10 (
	.BITSLIP((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed10),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[26]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[10]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[26]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[10]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[26]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[10]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[26]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[10])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_10 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay10),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed10)
);

IOBUF IOBUF_10(
	.I(soc_videosoc_ddrphy_dq_o10),
	.T(soc_videosoc_ddrphy_dq_t10),
	.IO(ddram_dq[10]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay10)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_40 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[11]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[27]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[11]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[27]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[11]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[27]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[11]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[27]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o11),
	.TQ(soc_videosoc_ddrphy_dq_t11)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_11 (
	.BITSLIP((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed11),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[27]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[11]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[27]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[11]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[27]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[11]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[27]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[11])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_11 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay11),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed11)
);

IOBUF IOBUF_11(
	.I(soc_videosoc_ddrphy_dq_o11),
	.T(soc_videosoc_ddrphy_dq_t11),
	.IO(ddram_dq[11]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay11)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_41 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[12]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[28]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[12]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[28]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[12]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[28]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[12]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[28]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o12),
	.TQ(soc_videosoc_ddrphy_dq_t12)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_12 (
	.BITSLIP((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed12),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[28]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[12]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[28]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[12]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[28]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[12]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[28]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[12])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_12 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay12),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed12)
);

IOBUF IOBUF_12(
	.I(soc_videosoc_ddrphy_dq_o12),
	.T(soc_videosoc_ddrphy_dq_t12),
	.IO(ddram_dq[12]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay12)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_42 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[13]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[29]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[13]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[29]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[13]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[29]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[13]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[29]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o13),
	.TQ(soc_videosoc_ddrphy_dq_t13)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_13 (
	.BITSLIP((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed13),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[29]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[13]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[29]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[13]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[29]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[13]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[29]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[13])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_13 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay13),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed13)
);

IOBUF IOBUF_13(
	.I(soc_videosoc_ddrphy_dq_o13),
	.T(soc_videosoc_ddrphy_dq_t13),
	.IO(ddram_dq[13]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay13)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_43 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[14]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[30]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[14]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[30]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[14]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[30]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[14]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[30]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o14),
	.TQ(soc_videosoc_ddrphy_dq_t14)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_14 (
	.BITSLIP((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed14),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[30]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[14]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[30]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[14]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[30]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[14]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[30]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[14])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_14 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay14),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed14)
);

IOBUF IOBUF_14(
	.I(soc_videosoc_ddrphy_dq_o14),
	.T(soc_videosoc_ddrphy_dq_t14),
	.IO(ddram_dq[14]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay14)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_44 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(soc_videosoc_ddrphy_dfi_p0_wrdata[15]),
	.D2(soc_videosoc_ddrphy_dfi_p0_wrdata[31]),
	.D3(soc_videosoc_ddrphy_dfi_p1_wrdata[15]),
	.D4(soc_videosoc_ddrphy_dfi_p1_wrdata[31]),
	.D5(soc_videosoc_ddrphy_dfi_p2_wrdata[15]),
	.D6(soc_videosoc_ddrphy_dfi_p2_wrdata[31]),
	.D7(soc_videosoc_ddrphy_dfi_p3_wrdata[15]),
	.D8(soc_videosoc_ddrphy_dfi_p3_wrdata[31]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~soc_videosoc_ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(soc_videosoc_ddrphy_dq_o15),
	.TQ(soc_videosoc_ddrphy_dq_t15)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_15 (
	.BITSLIP((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_bitslip_re)),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB((~sys4x_clk)),
	.CLKDIV(sys_clk),
	.DDLY(soc_videosoc_ddrphy_dq_i_delayed15),
	.RST((sys_rst | (soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re))),
	.Q1(soc_videosoc_ddrphy_dfi_p3_rddata[31]),
	.Q2(soc_videosoc_ddrphy_dfi_p3_rddata[15]),
	.Q3(soc_videosoc_ddrphy_dfi_p2_rddata[31]),
	.Q4(soc_videosoc_ddrphy_dfi_p2_rddata[15]),
	.Q5(soc_videosoc_ddrphy_dfi_p1_rddata[31]),
	.Q6(soc_videosoc_ddrphy_dfi_p1_rddata[15]),
	.Q7(soc_videosoc_ddrphy_dfi_p0_rddata[31]),
	.Q8(soc_videosoc_ddrphy_dfi_p0_rddata[15])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(3'd6),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_15 (
	.C(sys_clk),
	.CE((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_inc_re)),
	.IDATAIN(soc_videosoc_ddrphy_dq_i_nodelay15),
	.INC(1'd1),
	.LD((soc_videosoc_ddrphy_storage[1] & soc_videosoc_ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_videosoc_ddrphy_dq_i_delayed15)
);

IOBUF IOBUF_15(
	.I(soc_videosoc_ddrphy_dq_o15),
	.T(soc_videosoc_ddrphy_dq_t15),
	.IO(ddram_dq[15]),
	.O(soc_videosoc_ddrphy_dq_i_nodelay15)
);

reg [24:0] storage_2[0:7];
reg [2:0] memadr_3;
always @(posedge sys_clk) begin
	if (soc_videosoc_sdram_bankmachine0_wrport_we)
		storage_2[soc_videosoc_sdram_bankmachine0_wrport_adr] <= soc_videosoc_sdram_bankmachine0_wrport_dat_w;
	memadr_3 <= soc_videosoc_sdram_bankmachine0_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign soc_videosoc_sdram_bankmachine0_wrport_dat_r = storage_2[memadr_3];
assign soc_videosoc_sdram_bankmachine0_rdport_dat_r = storage_2[soc_videosoc_sdram_bankmachine0_rdport_adr];

reg [24:0] storage_3[0:7];
reg [2:0] memadr_4;
always @(posedge sys_clk) begin
	if (soc_videosoc_sdram_bankmachine1_wrport_we)
		storage_3[soc_videosoc_sdram_bankmachine1_wrport_adr] <= soc_videosoc_sdram_bankmachine1_wrport_dat_w;
	memadr_4 <= soc_videosoc_sdram_bankmachine1_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign soc_videosoc_sdram_bankmachine1_wrport_dat_r = storage_3[memadr_4];
assign soc_videosoc_sdram_bankmachine1_rdport_dat_r = storage_3[soc_videosoc_sdram_bankmachine1_rdport_adr];

reg [24:0] storage_4[0:7];
reg [2:0] memadr_5;
always @(posedge sys_clk) begin
	if (soc_videosoc_sdram_bankmachine2_wrport_we)
		storage_4[soc_videosoc_sdram_bankmachine2_wrport_adr] <= soc_videosoc_sdram_bankmachine2_wrport_dat_w;
	memadr_5 <= soc_videosoc_sdram_bankmachine2_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign soc_videosoc_sdram_bankmachine2_wrport_dat_r = storage_4[memadr_5];
assign soc_videosoc_sdram_bankmachine2_rdport_dat_r = storage_4[soc_videosoc_sdram_bankmachine2_rdport_adr];

reg [24:0] storage_5[0:7];
reg [2:0] memadr_6;
always @(posedge sys_clk) begin
	if (soc_videosoc_sdram_bankmachine3_wrport_we)
		storage_5[soc_videosoc_sdram_bankmachine3_wrport_adr] <= soc_videosoc_sdram_bankmachine3_wrport_dat_w;
	memadr_6 <= soc_videosoc_sdram_bankmachine3_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign soc_videosoc_sdram_bankmachine3_wrport_dat_r = storage_5[memadr_6];
assign soc_videosoc_sdram_bankmachine3_rdport_dat_r = storage_5[soc_videosoc_sdram_bankmachine3_rdport_adr];

reg [24:0] storage_6[0:7];
reg [2:0] memadr_7;
always @(posedge sys_clk) begin
	if (soc_videosoc_sdram_bankmachine4_wrport_we)
		storage_6[soc_videosoc_sdram_bankmachine4_wrport_adr] <= soc_videosoc_sdram_bankmachine4_wrport_dat_w;
	memadr_7 <= soc_videosoc_sdram_bankmachine4_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign soc_videosoc_sdram_bankmachine4_wrport_dat_r = storage_6[memadr_7];
assign soc_videosoc_sdram_bankmachine4_rdport_dat_r = storage_6[soc_videosoc_sdram_bankmachine4_rdport_adr];

reg [24:0] storage_7[0:7];
reg [2:0] memadr_8;
always @(posedge sys_clk) begin
	if (soc_videosoc_sdram_bankmachine5_wrport_we)
		storage_7[soc_videosoc_sdram_bankmachine5_wrport_adr] <= soc_videosoc_sdram_bankmachine5_wrport_dat_w;
	memadr_8 <= soc_videosoc_sdram_bankmachine5_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign soc_videosoc_sdram_bankmachine5_wrport_dat_r = storage_7[memadr_8];
assign soc_videosoc_sdram_bankmachine5_rdport_dat_r = storage_7[soc_videosoc_sdram_bankmachine5_rdport_adr];

reg [24:0] storage_8[0:7];
reg [2:0] memadr_9;
always @(posedge sys_clk) begin
	if (soc_videosoc_sdram_bankmachine6_wrport_we)
		storage_8[soc_videosoc_sdram_bankmachine6_wrport_adr] <= soc_videosoc_sdram_bankmachine6_wrport_dat_w;
	memadr_9 <= soc_videosoc_sdram_bankmachine6_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign soc_videosoc_sdram_bankmachine6_wrport_dat_r = storage_8[memadr_9];
assign soc_videosoc_sdram_bankmachine6_rdport_dat_r = storage_8[soc_videosoc_sdram_bankmachine6_rdport_adr];

reg [24:0] storage_9[0:7];
reg [2:0] memadr_10;
always @(posedge sys_clk) begin
	if (soc_videosoc_sdram_bankmachine7_wrport_we)
		storage_9[soc_videosoc_sdram_bankmachine7_wrport_adr] <= soc_videosoc_sdram_bankmachine7_wrport_dat_w;
	memadr_10 <= soc_videosoc_sdram_bankmachine7_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign soc_videosoc_sdram_bankmachine7_wrport_dat_r = storage_9[memadr_10];
assign soc_videosoc_sdram_bankmachine7_rdport_dat_r = storage_9[soc_videosoc_sdram_bankmachine7_rdport_adr];

reg [23:0] tag_mem[0:511];
reg [8:0] memadr_11;
always @(posedge sys_clk) begin
	if (soc_videosoc_tag_port_we)
		tag_mem[soc_videosoc_tag_port_adr] <= soc_videosoc_tag_port_dat_w;
	memadr_11 <= soc_videosoc_tag_port_adr;
end

assign soc_videosoc_tag_port_dat_r = tag_mem[memadr_11];

STARTUPE2 STARTUPE2(
	.CLK(1'd0),
	.GSR(1'd0),
	.GTS(1'd0),
	.KEYCLEARB(1'd0),
	.PACK(1'd0),
	.USRCCLKO(soc_videosoc_clk0),
	.USRCCLKTS(1'd0),
	.USRDONEO(1'd1),
	.USRDONETS(1'd1)
);

IBUF IBUF(
	.I(eth_clocks_rx),
	.O(soc_ethphy_eth_rx_clk_ibuf)
);

BUFG BUFG_5(
	.I(soc_ethphy_eth_rx_clk_ibuf),
	.O(eth_rx_clk)
);

PLLE2_BASE #(
	.CLKFBOUT_MULT(4'd8),
	.CLKIN1_PERIOD(8.0),
	.CLKOUT0_DIVIDE(4'd8),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(4'd8),
	.CLKOUT1_PHASE(90.0),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER1(0.01),
	.STARTUP_WAIT("FALSE")
) PLLE2_BASE_1 (
	.CLKFBIN(soc_ethphy_pll_fb),
	.CLKIN1(eth_rx_clk),
	.CLKFBOUT(soc_ethphy_pll_fb),
	.CLKOUT0(soc_ethphy_pll_clk_tx),
	.CLKOUT1(soc_ethphy_pll_clk_tx90),
	.LOCKED(soc_ethphy_pll_locked)
);

BUFG BUFG_6(
	.I(soc_ethphy_pll_clk_tx),
	.O(eth_tx_clk)
);

BUFG BUFG_7(
	.I(soc_ethphy_pll_clk_tx90),
	.O(eth_tx90_clk)
);

ODDR #(
	.DDR_CLK_EDGE("SAME_EDGE")
) ODDR (
	.C(eth_tx90_clk),
	.CE(1'd1),
	.D1(1'd1),
	.D2(1'd0),
	.R(1'd0),
	.S(1'd0),
	.Q(soc_ethphy_eth_tx_clk_obuf)
);

OBUF OBUF(
	.I(soc_ethphy_eth_tx_clk_obuf),
	.O(eth_clocks_tx)
);

ODDR #(
	.DDR_CLK_EDGE("SAME_EDGE")
) ODDR_1 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D1(soc_ethphy_sink_valid),
	.D2(soc_ethphy_sink_valid),
	.R(1'd0),
	.S(1'd0),
	.Q(soc_ethphy_tx_ctl_obuf)
);

OBUF OBUF_1(
	.I(soc_ethphy_tx_ctl_obuf),
	.O(eth_tx_ctl)
);

ODDR #(
	.DDR_CLK_EDGE("SAME_EDGE")
) ODDR_2 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D1(soc_ethphy_sink_payload_data[0]),
	.D2(soc_ethphy_sink_payload_data[4]),
	.R(1'd0),
	.S(1'd0),
	.Q(soc_ethphy_tx_data_obuf[0])
);

OBUF OBUF_2(
	.I(soc_ethphy_tx_data_obuf[0]),
	.O(eth_tx_data[0])
);

ODDR #(
	.DDR_CLK_EDGE("SAME_EDGE")
) ODDR_3 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D1(soc_ethphy_sink_payload_data[1]),
	.D2(soc_ethphy_sink_payload_data[5]),
	.R(1'd0),
	.S(1'd0),
	.Q(soc_ethphy_tx_data_obuf[1])
);

OBUF OBUF_3(
	.I(soc_ethphy_tx_data_obuf[1]),
	.O(eth_tx_data[1])
);

ODDR #(
	.DDR_CLK_EDGE("SAME_EDGE")
) ODDR_4 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D1(soc_ethphy_sink_payload_data[2]),
	.D2(soc_ethphy_sink_payload_data[6]),
	.R(1'd0),
	.S(1'd0),
	.Q(soc_ethphy_tx_data_obuf[2])
);

OBUF OBUF_4(
	.I(soc_ethphy_tx_data_obuf[2]),
	.O(eth_tx_data[2])
);

ODDR #(
	.DDR_CLK_EDGE("SAME_EDGE")
) ODDR_5 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D1(soc_ethphy_sink_payload_data[3]),
	.D2(soc_ethphy_sink_payload_data[7]),
	.R(1'd0),
	.S(1'd0),
	.Q(soc_ethphy_tx_data_obuf[3])
);

OBUF OBUF_5(
	.I(soc_ethphy_tx_data_obuf[3]),
	.O(eth_tx_data[3])
);

IBUF IBUF_1(
	.I(eth_rx_ctl),
	.O(soc_ethphy_rx_ctl_ibuf)
);

IDELAYE2 #(
	.IDELAY_TYPE("FIXED")
) IDELAYE2_16 (
	.C(1'd0),
	.CE(1'd0),
	.IDATAIN(soc_ethphy_rx_ctl_ibuf),
	.INC(1'd0),
	.LD(1'd0),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_ethphy_rx_ctl_idelay)
);

IDDR #(
	.DDR_CLK_EDGE("SAME_EDGE_PIPELINED")
) IDDR (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(soc_ethphy_rx_ctl_idelay),
	.R(1'd0),
	.S(1'd0),
	.Q1(soc_ethphy_rx_ctl)
);

IBUF IBUF_2(
	.I(eth_rx_data[0]),
	.O(soc_ethphy_rx_data_ibuf[0])
);

IDELAYE2 #(
	.IDELAY_TYPE("FIXED")
) IDELAYE2_17 (
	.C(1'd0),
	.CE(1'd0),
	.IDATAIN(soc_ethphy_rx_data_ibuf[0]),
	.INC(1'd0),
	.LD(1'd0),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_ethphy_rx_data_idelay[0])
);

IDDR #(
	.DDR_CLK_EDGE("SAME_EDGE_PIPELINED")
) IDDR_1 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(soc_ethphy_rx_data_idelay[0]),
	.R(1'd0),
	.S(1'd0),
	.Q1(soc_ethphy_rx_data[0]),
	.Q2(soc_ethphy_rx_data[4])
);

IBUF IBUF_3(
	.I(eth_rx_data[1]),
	.O(soc_ethphy_rx_data_ibuf[1])
);

IDELAYE2 #(
	.IDELAY_TYPE("FIXED")
) IDELAYE2_18 (
	.C(1'd0),
	.CE(1'd0),
	.IDATAIN(soc_ethphy_rx_data_ibuf[1]),
	.INC(1'd0),
	.LD(1'd0),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_ethphy_rx_data_idelay[1])
);

IDDR #(
	.DDR_CLK_EDGE("SAME_EDGE_PIPELINED")
) IDDR_2 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(soc_ethphy_rx_data_idelay[1]),
	.R(1'd0),
	.S(1'd0),
	.Q1(soc_ethphy_rx_data[1]),
	.Q2(soc_ethphy_rx_data[5])
);

IBUF IBUF_4(
	.I(eth_rx_data[2]),
	.O(soc_ethphy_rx_data_ibuf[2])
);

IDELAYE2 #(
	.IDELAY_TYPE("FIXED")
) IDELAYE2_19 (
	.C(1'd0),
	.CE(1'd0),
	.IDATAIN(soc_ethphy_rx_data_ibuf[2]),
	.INC(1'd0),
	.LD(1'd0),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_ethphy_rx_data_idelay[2])
);

IDDR #(
	.DDR_CLK_EDGE("SAME_EDGE_PIPELINED")
) IDDR_3 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(soc_ethphy_rx_data_idelay[2]),
	.R(1'd0),
	.S(1'd0),
	.Q1(soc_ethphy_rx_data[2]),
	.Q2(soc_ethphy_rx_data[6])
);

IBUF IBUF_5(
	.I(eth_rx_data[3]),
	.O(soc_ethphy_rx_data_ibuf[3])
);

IDELAYE2 #(
	.IDELAY_TYPE("FIXED")
) IDELAYE2_20 (
	.C(1'd0),
	.CE(1'd0),
	.IDATAIN(soc_ethphy_rx_data_ibuf[3]),
	.INC(1'd0),
	.LD(1'd0),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_ethphy_rx_data_idelay[3])
);

IDDR #(
	.DDR_CLK_EDGE("SAME_EDGE_PIPELINED")
) IDDR_4 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(soc_ethphy_rx_data_idelay[3]),
	.R(1'd0),
	.S(1'd0),
	.Q1(soc_ethphy_rx_data[3]),
	.Q2(soc_ethphy_rx_data[7])
);

assign eth_mdio = soc_ethphy_data_oe ? soc_ethphy_data_w : 1'bz;
assign soc_ethphy_data_r = eth_mdio;

reg [11:0] storage_10[0:4];
reg [2:0] memadr_12;
always @(posedge eth_rx_clk) begin
	if (soc_ethmac_crc32_checker_syncfifo_wrport_we)
		storage_10[soc_ethmac_crc32_checker_syncfifo_wrport_adr] <= soc_ethmac_crc32_checker_syncfifo_wrport_dat_w;
	memadr_12 <= soc_ethmac_crc32_checker_syncfifo_wrport_adr;
end

always @(posedge eth_rx_clk) begin
end

assign soc_ethmac_crc32_checker_syncfifo_wrport_dat_r = storage_10[memadr_12];
assign soc_ethmac_crc32_checker_syncfifo_rdport_dat_r = storage_10[soc_ethmac_crc32_checker_syncfifo_rdport_adr];

reg [41:0] storage_11[0:63];
reg [5:0] memadr_13;
reg [41:0] memdat_1;
always @(posedge sys_clk) begin
	if (soc_ethmac_tx_cdc_wrport_we)
		storage_11[soc_ethmac_tx_cdc_wrport_adr] <= soc_ethmac_tx_cdc_wrport_dat_w;
	memadr_13 <= soc_ethmac_tx_cdc_wrport_adr;
end

always @(posedge eth_tx_clk) begin
	memdat_1 <= storage_11[soc_ethmac_tx_cdc_rdport_adr];
end

assign soc_ethmac_tx_cdc_wrport_dat_r = storage_11[memadr_13];
assign soc_ethmac_tx_cdc_rdport_dat_r = memdat_1;

reg [41:0] storage_12[0:63];
reg [5:0] memadr_14;
reg [41:0] memdat_2;
always @(posedge eth_rx_clk) begin
	if (soc_ethmac_rx_cdc_wrport_we)
		storage_12[soc_ethmac_rx_cdc_wrport_adr] <= soc_ethmac_rx_cdc_wrport_dat_w;
	memadr_14 <= soc_ethmac_rx_cdc_wrport_adr;
end

always @(posedge sys_clk) begin
	memdat_2 <= storage_12[soc_ethmac_rx_cdc_rdport_adr];
end

assign soc_ethmac_rx_cdc_wrport_dat_r = storage_12[memadr_14];
assign soc_ethmac_rx_cdc_rdport_dat_r = memdat_2;

reg [34:0] storage_13[0:1];
reg [0:0] memadr_15;
always @(posedge sys_clk) begin
	if (soc_ethmac_writer_fifo_wrport_we)
		storage_13[soc_ethmac_writer_fifo_wrport_adr] <= soc_ethmac_writer_fifo_wrport_dat_w;
	memadr_15 <= soc_ethmac_writer_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign soc_ethmac_writer_fifo_wrport_dat_r = storage_13[memadr_15];
assign soc_ethmac_writer_fifo_rdport_dat_r = storage_13[soc_ethmac_writer_fifo_rdport_adr];

reg [31:0] mem_2[0:511];
reg [8:0] memadr_16;
reg [31:0] memdat_3;
always @(posedge sys_clk) begin
	if (soc_ethmac_writer_memory0_we)
		mem_2[soc_ethmac_writer_memory0_adr] <= soc_ethmac_writer_memory0_dat_w;
	memadr_16 <= soc_ethmac_writer_memory0_adr;
end

always @(posedge sys_clk) begin
	memdat_3 <= mem_2[soc_ethmac_sram0_adr0];
end

assign soc_ethmac_writer_memory0_dat_r = mem_2[memadr_16];
assign soc_ethmac_sram0_dat_r0 = memdat_3;

reg [31:0] mem_3[0:511];
reg [8:0] memadr_17;
reg [31:0] memdat_4;
always @(posedge sys_clk) begin
	if (soc_ethmac_writer_memory1_we)
		mem_3[soc_ethmac_writer_memory1_adr] <= soc_ethmac_writer_memory1_dat_w;
	memadr_17 <= soc_ethmac_writer_memory1_adr;
end

always @(posedge sys_clk) begin
	memdat_4 <= mem_3[soc_ethmac_sram1_adr0];
end

assign soc_ethmac_writer_memory1_dat_r = mem_3[memadr_17];
assign soc_ethmac_sram1_dat_r0 = memdat_4;

reg [13:0] storage_14[0:1];
reg [0:0] memadr_18;
always @(posedge sys_clk) begin
	if (soc_ethmac_reader_fifo_wrport_we)
		storage_14[soc_ethmac_reader_fifo_wrport_adr] <= soc_ethmac_reader_fifo_wrport_dat_w;
	memadr_18 <= soc_ethmac_reader_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign soc_ethmac_reader_fifo_wrport_dat_r = storage_14[memadr_18];
assign soc_ethmac_reader_fifo_rdport_dat_r = storage_14[soc_ethmac_reader_fifo_rdport_adr];

reg [7:0] edid_mem[0:127];
reg [7:0] memdat_5;
reg [6:0] memadr_19;
always @(posedge sys_clk) begin
	memdat_5 <= edid_mem[soc_edid_adr];
end

always @(posedge sys_clk) begin
	if (vns_videosoc_we)
		edid_mem[vns_videosoc_adr] <= vns_videosoc_dat_w;
	memadr_19 <= vns_videosoc_adr;
end

assign soc_edid_dat_r = memdat_5;
assign vns_videosoc_dat_r = edid_mem[memadr_19];

initial begin
	$readmemh("edid_mem.init", edid_mem);
end

assign hdmi_in_sda = soc_edid_sda_drv_reg ? 1'd0 : 1'bz;
assign soc_edid_sda_i_async = hdmi_in_sda;

IBUFDS hdmi_in_ibufds(
	.I(hdmi_in_clk_p),
	.IB(hdmi_in_clk_n),
	.O(soc_clk_input)
);

BUFG BUFG_8(
	.I(soc_clk_input),
	.O(soc_clk_input_bufg)
);

MMCME2_ADV #(
	.BANDWIDTH("OPTIMIZED"),
	.CLKFBOUT_MULT_F(10.0),
	.CLKFBOUT_PHASE(0.0),
	.CLKIN1_PERIOD(6.734006734006734),
	.CLKOUT0_DIVIDE_F(4'd10),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(4'd8),
	.CLKOUT1_PHASE(0.0),
	.CLKOUT2_DIVIDE(2'd2),
	.CLKOUT2_PHASE(0.0),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER1(0.01)
) MMCME2_ADV (
	.CLKFBIN(soc_mmcm_fb),
	.CLKIN1(soc_clk_input),
	.DADDR(soc_mmcm_adr_storage),
	.DCLK(sys_clk),
	.DEN((soc_mmcm_read_re | soc_mmcm_write_re)),
	.DI(soc_mmcm_dat_w_storage),
	.DWE(soc_mmcm_write_re),
	.RST(soc_mmcm_reset_storage),
	.CLKFBOUT(soc_mmcm_fb),
	.CLKOUT0(soc_mmcm_clk0),
	.CLKOUT1(soc_mmcm_clk1),
	.CLKOUT2(soc_mmcm_clk2),
	.DO(soc_mmcm_dat_r_status),
	.DRDY(soc_mmcm_drdy),
	.LOCKED(soc_mmcm_locked)
);

BUFG BUFG_9(
	.I(soc_mmcm_clk0),
	.O(hdmi_in0_pix_clk)
);

BUFR BUFR(
	.I(soc_mmcm_clk1),
	.O(pix1p25x_clk)
);

BUFIO BUFIO(
	.I(soc_mmcm_clk2),
	.O(hdmi_in0_pix5x_clk)
);

IBUFDS_DIFF_OUT IBUFDS_DIFF_OUT(
	.I(hdmi_in_data0_p),
	.IB(hdmi_in_data0_n),
	.O(soc_s7datacapture0_serdes_m_i_nodelay),
	.OB(soc_s7datacapture0_serdes_s_i_nodelay)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_21 (
	.C(pix1p25x_clk),
	.CE(soc_s7datacapture0_delay_master_ce),
	.IDATAIN(soc_s7datacapture0_serdes_m_i_nodelay),
	.INC(soc_s7datacapture0_delay_master_inc),
	.LD(soc_s7datacapture0_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_s7datacapture0_serdes_m_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_16 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(pix1p25x_clk),
	.DDLY(soc_s7datacapture0_serdes_m_i_delayed),
	.RST(pix1p25x_rst),
	.Q1(soc_s7datacapture0_serdes_m_q[7]),
	.Q2(soc_s7datacapture0_serdes_m_q[6]),
	.Q3(soc_s7datacapture0_serdes_m_q[5]),
	.Q4(soc_s7datacapture0_serdes_m_q[4]),
	.Q5(soc_s7datacapture0_serdes_m_q[3]),
	.Q6(soc_s7datacapture0_serdes_m_q[2]),
	.Q7(soc_s7datacapture0_serdes_m_q[1]),
	.Q8(soc_s7datacapture0_serdes_m_q[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_22 (
	.C(pix1p25x_clk),
	.CE(soc_s7datacapture0_delay_slave_ce),
	.IDATAIN(soc_s7datacapture0_serdes_s_i_nodelay),
	.INC(soc_s7datacapture0_delay_slave_inc),
	.LD(soc_s7datacapture0_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_s7datacapture0_serdes_s_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_17 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(pix1p25x_clk),
	.DDLY(soc_s7datacapture0_serdes_s_i_delayed),
	.RST(pix1p25x_rst),
	.Q1(soc_s7datacapture0_serdes_s_q[7]),
	.Q2(soc_s7datacapture0_serdes_s_q[6]),
	.Q3(soc_s7datacapture0_serdes_s_q[5]),
	.Q4(soc_s7datacapture0_serdes_s_q[4]),
	.Q5(soc_s7datacapture0_serdes_s_q[3]),
	.Q6(soc_s7datacapture0_serdes_s_q[2]),
	.Q7(soc_s7datacapture0_serdes_s_q[1]),
	.Q8(soc_s7datacapture0_serdes_s_q[0])
);

IBUFDS_DIFF_OUT IBUFDS_DIFF_OUT_1(
	.I(hdmi_in_data1_p),
	.IB(hdmi_in_data1_n),
	.O(soc_s7datacapture1_serdes_m_i_nodelay),
	.OB(soc_s7datacapture1_serdes_s_i_nodelay)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_23 (
	.C(pix1p25x_clk),
	.CE(soc_s7datacapture1_delay_master_ce),
	.IDATAIN(soc_s7datacapture1_serdes_m_i_nodelay),
	.INC(soc_s7datacapture1_delay_master_inc),
	.LD(soc_s7datacapture1_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_s7datacapture1_serdes_m_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_18 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(pix1p25x_clk),
	.DDLY(soc_s7datacapture1_serdes_m_i_delayed),
	.RST(pix1p25x_rst),
	.Q1(soc_s7datacapture1_serdes_m_q[7]),
	.Q2(soc_s7datacapture1_serdes_m_q[6]),
	.Q3(soc_s7datacapture1_serdes_m_q[5]),
	.Q4(soc_s7datacapture1_serdes_m_q[4]),
	.Q5(soc_s7datacapture1_serdes_m_q[3]),
	.Q6(soc_s7datacapture1_serdes_m_q[2]),
	.Q7(soc_s7datacapture1_serdes_m_q[1]),
	.Q8(soc_s7datacapture1_serdes_m_q[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_24 (
	.C(pix1p25x_clk),
	.CE(soc_s7datacapture1_delay_slave_ce),
	.IDATAIN(soc_s7datacapture1_serdes_s_i_nodelay),
	.INC(soc_s7datacapture1_delay_slave_inc),
	.LD(soc_s7datacapture1_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_s7datacapture1_serdes_s_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_19 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(pix1p25x_clk),
	.DDLY(soc_s7datacapture1_serdes_s_i_delayed),
	.RST(pix1p25x_rst),
	.Q1(soc_s7datacapture1_serdes_s_q[7]),
	.Q2(soc_s7datacapture1_serdes_s_q[6]),
	.Q3(soc_s7datacapture1_serdes_s_q[5]),
	.Q4(soc_s7datacapture1_serdes_s_q[4]),
	.Q5(soc_s7datacapture1_serdes_s_q[3]),
	.Q6(soc_s7datacapture1_serdes_s_q[2]),
	.Q7(soc_s7datacapture1_serdes_s_q[1]),
	.Q8(soc_s7datacapture1_serdes_s_q[0])
);

IBUFDS_DIFF_OUT IBUFDS_DIFF_OUT_2(
	.I(hdmi_in_data2_p),
	.IB(hdmi_in_data2_n),
	.O(soc_s7datacapture2_serdes_m_i_nodelay),
	.OB(soc_s7datacapture2_serdes_s_i_nodelay)
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_25 (
	.C(pix1p25x_clk),
	.CE(soc_s7datacapture2_delay_master_ce),
	.IDATAIN(soc_s7datacapture2_serdes_m_i_nodelay),
	.INC(soc_s7datacapture2_delay_master_inc),
	.LD(soc_s7datacapture2_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_s7datacapture2_serdes_m_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_20 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(pix1p25x_clk),
	.DDLY(soc_s7datacapture2_serdes_m_i_delayed),
	.RST(pix1p25x_rst),
	.Q1(soc_s7datacapture2_serdes_m_q[7]),
	.Q2(soc_s7datacapture2_serdes_m_q[6]),
	.Q3(soc_s7datacapture2_serdes_m_q[5]),
	.Q4(soc_s7datacapture2_serdes_m_q[4]),
	.Q5(soc_s7datacapture2_serdes_m_q[3]),
	.Q6(soc_s7datacapture2_serdes_m_q[2]),
	.Q7(soc_s7datacapture2_serdes_m_q[1]),
	.Q8(soc_s7datacapture2_serdes_m_q[0])
);

IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_26 (
	.C(pix1p25x_clk),
	.CE(soc_s7datacapture2_delay_slave_ce),
	.IDATAIN(soc_s7datacapture2_serdes_s_i_nodelay),
	.INC(soc_s7datacapture2_delay_slave_inc),
	.LD(soc_s7datacapture2_delay_rst),
	.LDPIPEEN(1'd0),
	.DATAOUT(soc_s7datacapture2_serdes_s_i_delayed)
);

ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_21 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(hdmi_in0_pix5x_clk),
	.CLKB((~hdmi_in0_pix5x_clk)),
	.CLKDIV(pix1p25x_clk),
	.DDLY(soc_s7datacapture2_serdes_s_i_delayed),
	.RST(pix1p25x_rst),
	.Q1(soc_s7datacapture2_serdes_s_q[7]),
	.Q2(soc_s7datacapture2_serdes_s_q[6]),
	.Q3(soc_s7datacapture2_serdes_s_q[5]),
	.Q4(soc_s7datacapture2_serdes_s_q[4]),
	.Q5(soc_s7datacapture2_serdes_s_q[3]),
	.Q6(soc_s7datacapture2_serdes_s_q[2]),
	.Q7(soc_s7datacapture2_serdes_s_q[1]),
	.Q8(soc_s7datacapture2_serdes_s_q[0])
);

reg [10:0] storage_15[0:7];
reg [2:0] memadr_20;
always @(posedge hdmi_in0_pix_clk) begin
	if (soc_chansync_syncbuffer0_wrport_we)
		storage_15[soc_chansync_syncbuffer0_wrport_adr] <= soc_chansync_syncbuffer0_wrport_dat_w;
	memadr_20 <= soc_chansync_syncbuffer0_wrport_adr;
end

always @(posedge hdmi_in0_pix_clk) begin
end

assign soc_chansync_syncbuffer0_wrport_dat_r = storage_15[memadr_20];
assign soc_chansync_syncbuffer0_rdport_dat_r = storage_15[soc_chansync_syncbuffer0_rdport_adr];

reg [10:0] storage_16[0:7];
reg [2:0] memadr_21;
always @(posedge hdmi_in0_pix_clk) begin
	if (soc_chansync_syncbuffer1_wrport_we)
		storage_16[soc_chansync_syncbuffer1_wrport_adr] <= soc_chansync_syncbuffer1_wrport_dat_w;
	memadr_21 <= soc_chansync_syncbuffer1_wrport_adr;
end

always @(posedge hdmi_in0_pix_clk) begin
end

assign soc_chansync_syncbuffer1_wrport_dat_r = storage_16[memadr_21];
assign soc_chansync_syncbuffer1_rdport_dat_r = storage_16[soc_chansync_syncbuffer1_rdport_adr];

reg [10:0] storage_17[0:7];
reg [2:0] memadr_22;
always @(posedge hdmi_in0_pix_clk) begin
	if (soc_chansync_syncbuffer2_wrport_we)
		storage_17[soc_chansync_syncbuffer2_wrport_adr] <= soc_chansync_syncbuffer2_wrport_dat_w;
	memadr_22 <= soc_chansync_syncbuffer2_wrport_adr;
end

always @(posedge hdmi_in0_pix_clk) begin
end

assign soc_chansync_syncbuffer2_wrport_dat_r = storage_17[memadr_22];
assign soc_chansync_syncbuffer2_rdport_dat_r = storage_17[soc_chansync_syncbuffer2_rdport_adr];

reg [130:0] storage_18[0:511];
reg [8:0] memadr_23;
reg [130:0] memdat_6;
always @(posedge hdmi_in0_pix_clk) begin
	if (soc_frame_fifo_wrport_we)
		storage_18[soc_frame_fifo_wrport_adr] <= soc_frame_fifo_wrport_dat_w;
	memadr_23 <= soc_frame_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
	memdat_6 <= storage_18[soc_frame_fifo_rdport_adr];
end

assign soc_frame_fifo_wrport_dat_r = storage_18[memadr_23];
assign soc_frame_fifo_rdport_dat_r = memdat_6;

reg [129:0] storage_19[0:15];
reg [3:0] memadr_24;
always @(posedge sys_clk) begin
	if (soc_dma_fifo_wrport_we)
		storage_19[soc_dma_fifo_wrport_adr] <= soc_dma_fifo_wrport_dat_w;
	memadr_24 <= soc_dma_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
end

assign soc_dma_fifo_wrport_dat_r = storage_19[memadr_24];
assign soc_dma_fifo_rdport_dat_r = storage_19[soc_dma_fifo_rdport_adr];

reg [27:0] storage_20[0:3];
reg [1:0] memadr_25;
reg [27:0] memdat_7;
always @(posedge hdmi_out0_pix_clk) begin
	if (soc_hdmi_out0_dram_port_cmd_fifo_wrport_we)
		storage_20[soc_hdmi_out0_dram_port_cmd_fifo_wrport_adr] <= soc_hdmi_out0_dram_port_cmd_fifo_wrport_dat_w;
	memadr_25 <= soc_hdmi_out0_dram_port_cmd_fifo_wrport_adr;
end

always @(posedge sys_clk) begin
	memdat_7 <= storage_20[soc_hdmi_out0_dram_port_cmd_fifo_rdport_adr];
end

assign soc_hdmi_out0_dram_port_cmd_fifo_wrport_dat_r = storage_20[memadr_25];
assign soc_hdmi_out0_dram_port_cmd_fifo_rdport_dat_r = memdat_7;

reg [129:0] storage_21[0:15];
reg [3:0] memadr_26;
reg [129:0] memdat_8;
always @(posedge sys_clk) begin
	if (soc_hdmi_out0_dram_port_rdata_fifo_wrport_we)
		storage_21[soc_hdmi_out0_dram_port_rdata_fifo_wrport_adr] <= soc_hdmi_out0_dram_port_rdata_fifo_wrport_dat_w;
	memadr_26 <= soc_hdmi_out0_dram_port_rdata_fifo_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
	memdat_8 <= storage_21[soc_hdmi_out0_dram_port_rdata_fifo_rdport_adr];
end

assign soc_hdmi_out0_dram_port_rdata_fifo_wrport_dat_r = storage_21[memadr_26];
assign soc_hdmi_out0_dram_port_rdata_fifo_rdport_dat_r = memdat_8;

reg [9:0] storage_22[0:3];
reg [1:0] memadr_27;
always @(posedge hdmi_out0_pix_clk) begin
	if (soc_hdmi_out0_dram_port_cmd_buffer_wrport_we)
		storage_22[soc_hdmi_out0_dram_port_cmd_buffer_wrport_adr] <= soc_hdmi_out0_dram_port_cmd_buffer_wrport_dat_w;
	memadr_27 <= soc_hdmi_out0_dram_port_cmd_buffer_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
end

assign soc_hdmi_out0_dram_port_cmd_buffer_wrport_dat_r = storage_22[memadr_27];
assign soc_hdmi_out0_dram_port_cmd_buffer_rdport_dat_r = storage_22[soc_hdmi_out0_dram_port_cmd_buffer_rdport_adr];

reg [161:0] storage_23[0:1];
reg [0:0] memadr_28;
reg [161:0] memdat_9;
always @(posedge sys_clk) begin
	if (soc_hdmi_out0_core_initiator_cdc_wrport_we)
		storage_23[soc_hdmi_out0_core_initiator_cdc_wrport_adr] <= soc_hdmi_out0_core_initiator_cdc_wrport_dat_w;
	memadr_28 <= soc_hdmi_out0_core_initiator_cdc_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
	memdat_9 <= storage_23[soc_hdmi_out0_core_initiator_cdc_rdport_adr];
end

assign soc_hdmi_out0_core_initiator_cdc_wrport_dat_r = storage_23[memadr_28];
assign soc_hdmi_out0_core_initiator_cdc_rdport_dat_r = memdat_9;

reg [17:0] storage_24[0:4095];
reg [11:0] memadr_29;
reg [17:0] memdat_10;
always @(posedge hdmi_out0_pix_clk) begin
	if (soc_hdmi_out0_core_dmareader_fifo_wrport_we)
		storage_24[soc_hdmi_out0_core_dmareader_fifo_wrport_adr] <= soc_hdmi_out0_core_dmareader_fifo_wrport_dat_w;
	memadr_29 <= soc_hdmi_out0_core_dmareader_fifo_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
	if (soc_hdmi_out0_core_dmareader_fifo_rdport_re)
		memdat_10 <= storage_24[soc_hdmi_out0_core_dmareader_fifo_rdport_adr];
end

assign soc_hdmi_out0_core_dmareader_fifo_wrport_dat_r = storage_24[memadr_29];
assign soc_hdmi_out0_core_dmareader_fifo_rdport_dat_r = memdat_10;

MMCME2_ADV #(
	.BANDWIDTH("OPTIMIZED"),
	.CLKFBOUT_MULT_F(30.0),
	.CLKFBOUT_PHASE(0.0),
	.CLKIN1_PERIOD(10.0),
	.CLKOUT0_DIVIDE_F(10.0),
	.CLKOUT0_PHASE(0.0),
	.CLKOUT1_DIVIDE(2'd2),
	.CLKOUT1_PHASE(0.0),
	.DIVCLK_DIVIDE(2'd2),
	.REF_JITTER1(0.01)
) MMCME2_ADV_1 (
	.CLKFBIN(soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_fb),
	.CLKIN1(clk100_clk),
	.DADDR(soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_adr_storage),
	.DCLK(sys_clk),
	.DEN((soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_read_re | soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_write_re)),
	.DI(soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_w_storage),
	.DWE(soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_write_re),
	.RST(soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_reset_storage),
	.CLKFBOUT(soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_fb),
	.CLKOUT0(soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_clk0),
	.CLKOUT1(soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_clk1),
	.DO(soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_dat_r_status),
	.DRDY(soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_drdy),
	.LOCKED(soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_locked)
);

BUFG BUFG_10(
	.I(soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_clk0),
	.O(hdmi_out0_pix_clk)
);

BUFG BUFG_11(
	.I(soc_hdmi_out0_driver_s7hdmioutclocking_mmcm_clk1),
	.O(hdmi_out0_pix5x_clk)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_45 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(soc_hdmi_out0_driver_s7hdmioutclocking_data1[0]),
	.D2(soc_hdmi_out0_driver_s7hdmioutclocking_data1[1]),
	.D3(soc_hdmi_out0_driver_s7hdmioutclocking_data1[2]),
	.D4(soc_hdmi_out0_driver_s7hdmioutclocking_data1[3]),
	.D5(soc_hdmi_out0_driver_s7hdmioutclocking_data1[4]),
	.D6(soc_hdmi_out0_driver_s7hdmioutclocking_data1[5]),
	.D7(soc_hdmi_out0_driver_s7hdmioutclocking_data1[6]),
	.D8(soc_hdmi_out0_driver_s7hdmioutclocking_data1[7]),
	.OCE(soc_hdmi_out0_driver_s7hdmioutclocking_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(soc_hdmi_out0_driver_s7hdmioutclocking_shift[0]),
	.SHIFTIN2(soc_hdmi_out0_driver_s7hdmioutclocking_shift[1]),
	.TCE(1'd0),
	.OQ(soc_hdmi_out0_driver_s7hdmioutclocking_pad_se)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("SLAVE"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_46 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(1'd0),
	.D2(1'd0),
	.D3(soc_hdmi_out0_driver_s7hdmioutclocking_data1[8]),
	.D4(soc_hdmi_out0_driver_s7hdmioutclocking_data1[9]),
	.D5(1'd0),
	.D6(1'd0),
	.D7(1'd0),
	.D8(1'd0),
	.OCE(soc_hdmi_out0_driver_s7hdmioutclocking_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.TCE(1'd0),
	.SHIFTOUT1(soc_hdmi_out0_driver_s7hdmioutclocking_shift[0]),
	.SHIFTOUT2(soc_hdmi_out0_driver_s7hdmioutclocking_shift[1])
);

OBUFDS OBUFDS_1(
	.I(soc_hdmi_out0_driver_s7hdmioutclocking_pad_se),
	.O(hdmi_out_clk_p),
	.OB(hdmi_out_clk_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_47 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(soc_hdmi_out0_driver_hdmi_phy_es0_data[0]),
	.D2(soc_hdmi_out0_driver_hdmi_phy_es0_data[1]),
	.D3(soc_hdmi_out0_driver_hdmi_phy_es0_data[2]),
	.D4(soc_hdmi_out0_driver_hdmi_phy_es0_data[3]),
	.D5(soc_hdmi_out0_driver_hdmi_phy_es0_data[4]),
	.D6(soc_hdmi_out0_driver_hdmi_phy_es0_data[5]),
	.D7(soc_hdmi_out0_driver_hdmi_phy_es0_data[6]),
	.D8(soc_hdmi_out0_driver_hdmi_phy_es0_data[7]),
	.OCE(soc_hdmi_out0_driver_hdmi_phy_es0_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(soc_hdmi_out0_driver_hdmi_phy_es0_shift[0]),
	.SHIFTIN2(soc_hdmi_out0_driver_hdmi_phy_es0_shift[1]),
	.TCE(1'd0),
	.OQ(soc_hdmi_out0_driver_hdmi_phy_es0_pad_se)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("SLAVE"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_48 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(1'd0),
	.D2(1'd0),
	.D3(soc_hdmi_out0_driver_hdmi_phy_es0_data[8]),
	.D4(soc_hdmi_out0_driver_hdmi_phy_es0_data[9]),
	.D5(1'd0),
	.D6(1'd0),
	.D7(1'd0),
	.D8(1'd0),
	.OCE(soc_hdmi_out0_driver_hdmi_phy_es0_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.TCE(1'd0),
	.SHIFTOUT1(soc_hdmi_out0_driver_hdmi_phy_es0_shift[0]),
	.SHIFTOUT2(soc_hdmi_out0_driver_hdmi_phy_es0_shift[1])
);

OBUFDS OBUFDS_2(
	.I(soc_hdmi_out0_driver_hdmi_phy_es0_pad_se),
	.O(hdmi_out_data0_p),
	.OB(hdmi_out_data0_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_49 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(soc_hdmi_out0_driver_hdmi_phy_es1_data[0]),
	.D2(soc_hdmi_out0_driver_hdmi_phy_es1_data[1]),
	.D3(soc_hdmi_out0_driver_hdmi_phy_es1_data[2]),
	.D4(soc_hdmi_out0_driver_hdmi_phy_es1_data[3]),
	.D5(soc_hdmi_out0_driver_hdmi_phy_es1_data[4]),
	.D6(soc_hdmi_out0_driver_hdmi_phy_es1_data[5]),
	.D7(soc_hdmi_out0_driver_hdmi_phy_es1_data[6]),
	.D8(soc_hdmi_out0_driver_hdmi_phy_es1_data[7]),
	.OCE(soc_hdmi_out0_driver_hdmi_phy_es1_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(soc_hdmi_out0_driver_hdmi_phy_es1_shift[0]),
	.SHIFTIN2(soc_hdmi_out0_driver_hdmi_phy_es1_shift[1]),
	.TCE(1'd0),
	.OQ(soc_hdmi_out0_driver_hdmi_phy_es1_pad_se)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("SLAVE"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_50 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(1'd0),
	.D2(1'd0),
	.D3(soc_hdmi_out0_driver_hdmi_phy_es1_data[8]),
	.D4(soc_hdmi_out0_driver_hdmi_phy_es1_data[9]),
	.D5(1'd0),
	.D6(1'd0),
	.D7(1'd0),
	.D8(1'd0),
	.OCE(soc_hdmi_out0_driver_hdmi_phy_es1_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.TCE(1'd0),
	.SHIFTOUT1(soc_hdmi_out0_driver_hdmi_phy_es1_shift[0]),
	.SHIFTOUT2(soc_hdmi_out0_driver_hdmi_phy_es1_shift[1])
);

OBUFDS OBUFDS_3(
	.I(soc_hdmi_out0_driver_hdmi_phy_es1_pad_se),
	.O(hdmi_out_data1_p),
	.OB(hdmi_out_data1_n)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_51 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(soc_hdmi_out0_driver_hdmi_phy_es2_data[0]),
	.D2(soc_hdmi_out0_driver_hdmi_phy_es2_data[1]),
	.D3(soc_hdmi_out0_driver_hdmi_phy_es2_data[2]),
	.D4(soc_hdmi_out0_driver_hdmi_phy_es2_data[3]),
	.D5(soc_hdmi_out0_driver_hdmi_phy_es2_data[4]),
	.D6(soc_hdmi_out0_driver_hdmi_phy_es2_data[5]),
	.D7(soc_hdmi_out0_driver_hdmi_phy_es2_data[6]),
	.D8(soc_hdmi_out0_driver_hdmi_phy_es2_data[7]),
	.OCE(soc_hdmi_out0_driver_hdmi_phy_es2_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(soc_hdmi_out0_driver_hdmi_phy_es2_shift[0]),
	.SHIFTIN2(soc_hdmi_out0_driver_hdmi_phy_es2_shift[1]),
	.TCE(1'd0),
	.OQ(soc_hdmi_out0_driver_hdmi_phy_es2_pad_se)
);

OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("DDR"),
	.DATA_WIDTH(4'd10),
	.SERDES_MODE("SLAVE"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_52 (
	.CLK(hdmi_out0_pix5x_clk),
	.CLKDIV(hdmi_out0_pix_clk),
	.D1(1'd0),
	.D2(1'd0),
	.D3(soc_hdmi_out0_driver_hdmi_phy_es2_data[8]),
	.D4(soc_hdmi_out0_driver_hdmi_phy_es2_data[9]),
	.D5(1'd0),
	.D6(1'd0),
	.D7(1'd0),
	.D8(1'd0),
	.OCE(soc_hdmi_out0_driver_hdmi_phy_es2_ce),
	.RST(hdmi_out0_pix_rst),
	.SHIFTIN1(1'd0),
	.SHIFTIN2(1'd0),
	.TCE(1'd0),
	.SHIFTOUT1(soc_hdmi_out0_driver_hdmi_phy_es2_shift[0]),
	.SHIFTOUT2(soc_hdmi_out0_driver_hdmi_phy_es2_shift[1])
);

OBUFDS OBUFDS_4(
	.I(soc_hdmi_out0_driver_hdmi_phy_es2_pad_se),
	.O(hdmi_out_data2_p),
	.OB(hdmi_out_data2_n)
);

reg [9:0] storage_25[0:3];
reg [1:0] memadr_30;
always @(posedge hdmi_out0_pix_clk) begin
	if (soc_hdmi_out0_resetinserter_y_fifo_wrport_we)
		storage_25[soc_hdmi_out0_resetinserter_y_fifo_wrport_adr] <= soc_hdmi_out0_resetinserter_y_fifo_wrport_dat_w;
	memadr_30 <= soc_hdmi_out0_resetinserter_y_fifo_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
end

assign soc_hdmi_out0_resetinserter_y_fifo_wrport_dat_r = storage_25[memadr_30];
assign soc_hdmi_out0_resetinserter_y_fifo_rdport_dat_r = storage_25[soc_hdmi_out0_resetinserter_y_fifo_rdport_adr];

reg [9:0] storage_26[0:3];
reg [1:0] memadr_31;
always @(posedge hdmi_out0_pix_clk) begin
	if (soc_hdmi_out0_resetinserter_cb_fifo_wrport_we)
		storage_26[soc_hdmi_out0_resetinserter_cb_fifo_wrport_adr] <= soc_hdmi_out0_resetinserter_cb_fifo_wrport_dat_w;
	memadr_31 <= soc_hdmi_out0_resetinserter_cb_fifo_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
end

assign soc_hdmi_out0_resetinserter_cb_fifo_wrport_dat_r = storage_26[memadr_31];
assign soc_hdmi_out0_resetinserter_cb_fifo_rdport_dat_r = storage_26[soc_hdmi_out0_resetinserter_cb_fifo_rdport_adr];

reg [9:0] storage_27[0:3];
reg [1:0] memadr_32;
always @(posedge hdmi_out0_pix_clk) begin
	if (soc_hdmi_out0_resetinserter_cr_fifo_wrport_we)
		storage_27[soc_hdmi_out0_resetinserter_cr_fifo_wrport_adr] <= soc_hdmi_out0_resetinserter_cr_fifo_wrport_dat_w;
	memadr_32 <= soc_hdmi_out0_resetinserter_cr_fifo_wrport_adr;
end

always @(posedge hdmi_out0_pix_clk) begin
end

assign soc_hdmi_out0_resetinserter_cr_fifo_wrport_dat_r = storage_27[memadr_32];
assign soc_hdmi_out0_resetinserter_cr_fifo_rdport_dat_r = storage_27[soc_hdmi_out0_resetinserter_cr_fifo_rdport_adr];

reg [7:0] data_mem_grain0[0:511];
reg [8:0] memadr_33;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[0])
		data_mem_grain0[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[7:0];
	memadr_33 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[7:0] = data_mem_grain0[memadr_33];

reg [7:0] data_mem_grain1[0:511];
reg [8:0] memadr_34;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[1])
		data_mem_grain1[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[15:8];
	memadr_34 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[15:8] = data_mem_grain1[memadr_34];

reg [7:0] data_mem_grain2[0:511];
reg [8:0] memadr_35;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[2])
		data_mem_grain2[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[23:16];
	memadr_35 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[23:16] = data_mem_grain2[memadr_35];

reg [7:0] data_mem_grain3[0:511];
reg [8:0] memadr_36;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[3])
		data_mem_grain3[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[31:24];
	memadr_36 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[31:24] = data_mem_grain3[memadr_36];

reg [7:0] data_mem_grain4[0:511];
reg [8:0] memadr_37;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[4])
		data_mem_grain4[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[39:32];
	memadr_37 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[39:32] = data_mem_grain4[memadr_37];

reg [7:0] data_mem_grain5[0:511];
reg [8:0] memadr_38;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[5])
		data_mem_grain5[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[47:40];
	memadr_38 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[47:40] = data_mem_grain5[memadr_38];

reg [7:0] data_mem_grain6[0:511];
reg [8:0] memadr_39;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[6])
		data_mem_grain6[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[55:48];
	memadr_39 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[55:48] = data_mem_grain6[memadr_39];

reg [7:0] data_mem_grain7[0:511];
reg [8:0] memadr_40;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[7])
		data_mem_grain7[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[63:56];
	memadr_40 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[63:56] = data_mem_grain7[memadr_40];

reg [7:0] data_mem_grain8[0:511];
reg [8:0] memadr_41;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[8])
		data_mem_grain8[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[71:64];
	memadr_41 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[71:64] = data_mem_grain8[memadr_41];

reg [7:0] data_mem_grain9[0:511];
reg [8:0] memadr_42;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[9])
		data_mem_grain9[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[79:72];
	memadr_42 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[79:72] = data_mem_grain9[memadr_42];

reg [7:0] data_mem_grain10[0:511];
reg [8:0] memadr_43;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[10])
		data_mem_grain10[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[87:80];
	memadr_43 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[87:80] = data_mem_grain10[memadr_43];

reg [7:0] data_mem_grain11[0:511];
reg [8:0] memadr_44;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[11])
		data_mem_grain11[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[95:88];
	memadr_44 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[95:88] = data_mem_grain11[memadr_44];

reg [7:0] data_mem_grain12[0:511];
reg [8:0] memadr_45;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[12])
		data_mem_grain12[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[103:96];
	memadr_45 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[103:96] = data_mem_grain12[memadr_45];

reg [7:0] data_mem_grain13[0:511];
reg [8:0] memadr_46;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[13])
		data_mem_grain13[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[111:104];
	memadr_46 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[111:104] = data_mem_grain13[memadr_46];

reg [7:0] data_mem_grain14[0:511];
reg [8:0] memadr_47;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[14])
		data_mem_grain14[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[119:112];
	memadr_47 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[119:112] = data_mem_grain14[memadr_47];

reg [7:0] data_mem_grain15[0:511];
reg [8:0] memadr_48;
always @(posedge sys_clk) begin
	if (soc_videosoc_data_port_we[15])
		data_mem_grain15[soc_videosoc_data_port_adr] <= soc_videosoc_data_port_dat_w[127:120];
	memadr_48 <= soc_videosoc_data_port_adr;
end

assign soc_videosoc_data_port_dat_r[127:120] = data_mem_grain15[memadr_48];

reg [7:0] mem_grain0[0:511];
reg [7:0] memdat_11;
reg [8:0] memadr_49;
always @(posedge sys_clk) begin
	memdat_11 <= mem_grain0[soc_ethmac_reader_memory0_adr];
end

always @(posedge sys_clk) begin
	if (soc_ethmac_sram0_we[0])
		mem_grain0[soc_ethmac_sram0_adr1] <= soc_ethmac_sram0_dat_w[7:0];
	memadr_49 <= soc_ethmac_sram0_adr1;
end

assign soc_ethmac_reader_memory0_dat_r[7:0] = memdat_11;
assign soc_ethmac_sram0_dat_r1[7:0] = mem_grain0[memadr_49];

reg [7:0] mem_grain1[0:511];
reg [7:0] memdat_12;
reg [8:0] memadr_50;
always @(posedge sys_clk) begin
	memdat_12 <= mem_grain1[soc_ethmac_reader_memory0_adr];
end

always @(posedge sys_clk) begin
	if (soc_ethmac_sram0_we[1])
		mem_grain1[soc_ethmac_sram0_adr1] <= soc_ethmac_sram0_dat_w[15:8];
	memadr_50 <= soc_ethmac_sram0_adr1;
end

assign soc_ethmac_reader_memory0_dat_r[15:8] = memdat_12;
assign soc_ethmac_sram0_dat_r1[15:8] = mem_grain1[memadr_50];

reg [7:0] mem_grain2[0:511];
reg [7:0] memdat_13;
reg [8:0] memadr_51;
always @(posedge sys_clk) begin
	memdat_13 <= mem_grain2[soc_ethmac_reader_memory0_adr];
end

always @(posedge sys_clk) begin
	if (soc_ethmac_sram0_we[2])
		mem_grain2[soc_ethmac_sram0_adr1] <= soc_ethmac_sram0_dat_w[23:16];
	memadr_51 <= soc_ethmac_sram0_adr1;
end

assign soc_ethmac_reader_memory0_dat_r[23:16] = memdat_13;
assign soc_ethmac_sram0_dat_r1[23:16] = mem_grain2[memadr_51];

reg [7:0] mem_grain3[0:511];
reg [7:0] memdat_14;
reg [8:0] memadr_52;
always @(posedge sys_clk) begin
	memdat_14 <= mem_grain3[soc_ethmac_reader_memory0_adr];
end

always @(posedge sys_clk) begin
	if (soc_ethmac_sram0_we[3])
		mem_grain3[soc_ethmac_sram0_adr1] <= soc_ethmac_sram0_dat_w[31:24];
	memadr_52 <= soc_ethmac_sram0_adr1;
end

assign soc_ethmac_reader_memory0_dat_r[31:24] = memdat_14;
assign soc_ethmac_sram0_dat_r1[31:24] = mem_grain3[memadr_52];

reg [7:0] mem_grain0_1[0:511];
reg [7:0] memdat_15;
reg [8:0] memadr_53;
always @(posedge sys_clk) begin
	memdat_15 <= mem_grain0_1[soc_ethmac_reader_memory1_adr];
end

always @(posedge sys_clk) begin
	if (soc_ethmac_sram1_we[0])
		mem_grain0_1[soc_ethmac_sram1_adr1] <= soc_ethmac_sram1_dat_w[7:0];
	memadr_53 <= soc_ethmac_sram1_adr1;
end

assign soc_ethmac_reader_memory1_dat_r[7:0] = memdat_15;
assign soc_ethmac_sram1_dat_r1[7:0] = mem_grain0_1[memadr_53];

reg [7:0] mem_grain1_1[0:511];
reg [7:0] memdat_16;
reg [8:0] memadr_54;
always @(posedge sys_clk) begin
	memdat_16 <= mem_grain1_1[soc_ethmac_reader_memory1_adr];
end

always @(posedge sys_clk) begin
	if (soc_ethmac_sram1_we[1])
		mem_grain1_1[soc_ethmac_sram1_adr1] <= soc_ethmac_sram1_dat_w[15:8];
	memadr_54 <= soc_ethmac_sram1_adr1;
end

assign soc_ethmac_reader_memory1_dat_r[15:8] = memdat_16;
assign soc_ethmac_sram1_dat_r1[15:8] = mem_grain1_1[memadr_54];

reg [7:0] mem_grain2_1[0:511];
reg [7:0] memdat_17;
reg [8:0] memadr_55;
always @(posedge sys_clk) begin
	memdat_17 <= mem_grain2_1[soc_ethmac_reader_memory1_adr];
end

always @(posedge sys_clk) begin
	if (soc_ethmac_sram1_we[2])
		mem_grain2_1[soc_ethmac_sram1_adr1] <= soc_ethmac_sram1_dat_w[23:16];
	memadr_55 <= soc_ethmac_sram1_adr1;
end

assign soc_ethmac_reader_memory1_dat_r[23:16] = memdat_17;
assign soc_ethmac_sram1_dat_r1[23:16] = mem_grain2_1[memadr_55];

reg [7:0] mem_grain3_1[0:511];
reg [7:0] memdat_18;
reg [8:0] memadr_56;
always @(posedge sys_clk) begin
	memdat_18 <= mem_grain3_1[soc_ethmac_reader_memory1_adr];
end

always @(posedge sys_clk) begin
	if (soc_ethmac_sram1_we[3])
		mem_grain3_1[soc_ethmac_sram1_adr1] <= soc_ethmac_sram1_dat_w[31:24];
	memadr_56 <= soc_ethmac_sram1_adr1;
end

assign soc_ethmac_reader_memory1_dat_r[31:24] = memdat_18;
assign soc_ethmac_sram1_dat_r1[31:24] = mem_grain3_1[memadr_56];

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE (
	.C(sys_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(vns_xilinxasyncresetsynchronizerimpl0),
	.Q(vns_xilinxasyncresetsynchronizerimpl0_rst_meta)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_1 (
	.C(sys_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl0_rst_meta),
	.PRE(vns_xilinxasyncresetsynchronizerimpl0),
	.Q(sys_rst)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_2 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(vns_xilinxasyncresetsynchronizerimpl1),
	.Q(vns_xilinxasyncresetsynchronizerimpl1_rst_meta)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_3 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl1_rst_meta),
	.PRE(vns_xilinxasyncresetsynchronizerimpl1),
	.Q(clk200_rst)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_4 (
	.C(clk100_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(vns_xilinxasyncresetsynchronizerimpl2),
	.Q(vns_xilinxasyncresetsynchronizerimpl2_rst_meta)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_5 (
	.C(clk100_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl2_rst_meta),
	.PRE(vns_xilinxasyncresetsynchronizerimpl2),
	.Q(clk100_rst)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_6 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(soc_ethphy_reset0),
	.Q(vns_xilinxasyncresetsynchronizerimpl3_rst_meta)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_7 (
	.C(eth_tx_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl3_rst_meta),
	.PRE(soc_ethphy_reset0),
	.Q(eth_tx_rst)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_8 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(soc_ethphy_reset0),
	.Q(vns_xilinxasyncresetsynchronizerimpl4_rst_meta)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_9 (
	.C(eth_rx_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl4_rst_meta),
	.PRE(soc_ethphy_reset0),
	.Q(eth_rx_rst)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_10 (
	.C(hdmi_in0_pix_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(vns_xilinxasyncresetsynchronizerimpl5),
	.Q(vns_xilinxasyncresetsynchronizerimpl5_rst_meta)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_11 (
	.C(hdmi_in0_pix_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl5_rst_meta),
	.PRE(vns_xilinxasyncresetsynchronizerimpl5),
	.Q(hdmi_in0_pix_rst)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_12 (
	.C(pix1p25x_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(vns_xilinxasyncresetsynchronizerimpl6),
	.Q(vns_xilinxasyncresetsynchronizerimpl6_rst_meta)
);

(* ars_ff = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_13 (
	.C(pix1p25x_clk),
	.CE(1'd1),
	.D(vns_xilinxasyncresetsynchronizerimpl6_rst_meta),
	.PRE(vns_xilinxasyncresetsynchronizerimpl6),
	.Q(pix1p25x_rst)
);

endmodule
